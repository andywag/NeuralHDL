//-----------------------------------------------------------------------------
// Company: 			                                                              
// Author:				Andy                                                          
// Date:                                                                       
// Module Name:       neuronStage
// Description:                                                                
//                                                                             
//-----------------------------------------------------------------------------

`ifndef TYPES
  `include "types.v"
  `define TYPES
`endif

    module neuronStage(
  input float_24_8              biasIn_0,
  input                         clk,
  input float_24_8              dataIn_0,
  input                         reset,
  input float_24_8              tapIn_0,
  input float_24_8              tapIn_1,
  input float_24_8              tapIn_10,
  input float_24_8              tapIn_100,
  input float_24_8              tapIn_101,
  input float_24_8              tapIn_102,
  input float_24_8              tapIn_103,
  input float_24_8              tapIn_104,
  input float_24_8              tapIn_105,
  input float_24_8              tapIn_106,
  input float_24_8              tapIn_107,
  input float_24_8              tapIn_108,
  input float_24_8              tapIn_109,
  input float_24_8              tapIn_11,
  input float_24_8              tapIn_110,
  input float_24_8              tapIn_111,
  input float_24_8              tapIn_112,
  input float_24_8              tapIn_113,
  input float_24_8              tapIn_114,
  input float_24_8              tapIn_115,
  input float_24_8              tapIn_116,
  input float_24_8              tapIn_117,
  input float_24_8              tapIn_118,
  input float_24_8              tapIn_119,
  input float_24_8              tapIn_12,
  input float_24_8              tapIn_120,
  input float_24_8              tapIn_121,
  input float_24_8              tapIn_122,
  input float_24_8              tapIn_123,
  input float_24_8              tapIn_124,
  input float_24_8              tapIn_125,
  input float_24_8              tapIn_126,
  input float_24_8              tapIn_127,
  input float_24_8              tapIn_13,
  input float_24_8              tapIn_14,
  input float_24_8              tapIn_15,
  input float_24_8              tapIn_16,
  input float_24_8              tapIn_17,
  input float_24_8              tapIn_18,
  input float_24_8              tapIn_19,
  input float_24_8              tapIn_2,
  input float_24_8              tapIn_20,
  input float_24_8              tapIn_21,
  input float_24_8              tapIn_22,
  input float_24_8              tapIn_23,
  input float_24_8              tapIn_24,
  input float_24_8              tapIn_25,
  input float_24_8              tapIn_26,
  input float_24_8              tapIn_27,
  input float_24_8              tapIn_28,
  input float_24_8              tapIn_29,
  input float_24_8              tapIn_3,
  input float_24_8              tapIn_30,
  input float_24_8              tapIn_31,
  input float_24_8              tapIn_32,
  input float_24_8              tapIn_33,
  input float_24_8              tapIn_34,
  input float_24_8              tapIn_35,
  input float_24_8              tapIn_36,
  input float_24_8              tapIn_37,
  input float_24_8              tapIn_38,
  input float_24_8              tapIn_39,
  input float_24_8              tapIn_4,
  input float_24_8              tapIn_40,
  input float_24_8              tapIn_41,
  input float_24_8              tapIn_42,
  input float_24_8              tapIn_43,
  input float_24_8              tapIn_44,
  input float_24_8              tapIn_45,
  input float_24_8              tapIn_46,
  input float_24_8              tapIn_47,
  input float_24_8              tapIn_48,
  input float_24_8              tapIn_49,
  input float_24_8              tapIn_5,
  input float_24_8              tapIn_50,
  input float_24_8              tapIn_51,
  input float_24_8              tapIn_52,
  input float_24_8              tapIn_53,
  input float_24_8              tapIn_54,
  input float_24_8              tapIn_55,
  input float_24_8              tapIn_56,
  input float_24_8              tapIn_57,
  input float_24_8              tapIn_58,
  input float_24_8              tapIn_59,
  input float_24_8              tapIn_6,
  input float_24_8              tapIn_60,
  input float_24_8              tapIn_61,
  input float_24_8              tapIn_62,
  input float_24_8              tapIn_63,
  input float_24_8              tapIn_64,
  input float_24_8              tapIn_65,
  input float_24_8              tapIn_66,
  input float_24_8              tapIn_67,
  input float_24_8              tapIn_68,
  input float_24_8              tapIn_69,
  input float_24_8              tapIn_7,
  input float_24_8              tapIn_70,
  input float_24_8              tapIn_71,
  input float_24_8              tapIn_72,
  input float_24_8              tapIn_73,
  input float_24_8              tapIn_74,
  input float_24_8              tapIn_75,
  input float_24_8              tapIn_76,
  input float_24_8              tapIn_77,
  input float_24_8              tapIn_78,
  input float_24_8              tapIn_79,
  input float_24_8              tapIn_8,
  input float_24_8              tapIn_80,
  input float_24_8              tapIn_81,
  input float_24_8              tapIn_82,
  input float_24_8              tapIn_83,
  input float_24_8              tapIn_84,
  input float_24_8              tapIn_85,
  input float_24_8              tapIn_86,
  input float_24_8              tapIn_87,
  input float_24_8              tapIn_88,
  input float_24_8              tapIn_89,
  input float_24_8              tapIn_9,
  input float_24_8              tapIn_90,
  input float_24_8              tapIn_91,
  input float_24_8              tapIn_92,
  input float_24_8              tapIn_93,
  input float_24_8              tapIn_94,
  input float_24_8              tapIn_95,
  input float_24_8              tapIn_96,
  input float_24_8              tapIn_97,
  input float_24_8              tapIn_98,
  input float_24_8              tapIn_99,
  input                         valid,
  output float_24_8             dataOutPre_0,
  output float_24_8             dataOut_0);

// Parameters 



// Wires 

  float_24_8                    biasIn_0_w0;  // <1,0>
  float_24_8                    biasIn_0_w1;  // <1,0>
  float_24_8                    biasIn_0_w10;  // <1,0>
  float_24_8                    biasIn_0_w100;  // <1,0>
  float_24_8                    biasIn_0_w101;  // <1,0>
  float_24_8                    biasIn_0_w102;  // <1,0>
  float_24_8                    biasIn_0_w103;  // <1,0>
  float_24_8                    biasIn_0_w104;  // <1,0>
  float_24_8                    biasIn_0_w105;  // <1,0>
  float_24_8                    biasIn_0_w106;  // <1,0>
  float_24_8                    biasIn_0_w107;  // <1,0>
  float_24_8                    biasIn_0_w108;  // <1,0>
  float_24_8                    biasIn_0_w109;  // <1,0>
  float_24_8                    biasIn_0_w11;  // <1,0>
  float_24_8                    biasIn_0_w110;  // <1,0>
  float_24_8                    biasIn_0_w111;  // <1,0>
  float_24_8                    biasIn_0_w112;  // <1,0>
  float_24_8                    biasIn_0_w113;  // <1,0>
  float_24_8                    biasIn_0_w114;  // <1,0>
  float_24_8                    biasIn_0_w115;  // <1,0>
  float_24_8                    biasIn_0_w116;  // <1,0>
  float_24_8                    biasIn_0_w117;  // <1,0>
  float_24_8                    biasIn_0_w118;  // <1,0>
  float_24_8                    biasIn_0_w119;  // <1,0>
  float_24_8                    biasIn_0_w12;  // <1,0>
  float_24_8                    biasIn_0_w120;  // <1,0>
  float_24_8                    biasIn_0_w121;  // <1,0>
  float_24_8                    biasIn_0_w122;  // <1,0>
  float_24_8                    biasIn_0_w123;  // <1,0>
  float_24_8                    biasIn_0_w124;  // <1,0>
  float_24_8                    biasIn_0_w125;  // <1,0>
  float_24_8                    biasIn_0_w126;  // <1,0>
  float_24_8                    biasIn_0_w127;  // <1,0>
  float_24_8                    biasIn_0_w13;  // <1,0>
  float_24_8                    biasIn_0_w14;  // <1,0>
  float_24_8                    biasIn_0_w15;  // <1,0>
  float_24_8                    biasIn_0_w16;  // <1,0>
  float_24_8                    biasIn_0_w17;  // <1,0>
  float_24_8                    biasIn_0_w18;  // <1,0>
  float_24_8                    biasIn_0_w19;  // <1,0>
  float_24_8                    biasIn_0_w2;  // <1,0>
  float_24_8                    biasIn_0_w20;  // <1,0>
  float_24_8                    biasIn_0_w21;  // <1,0>
  float_24_8                    biasIn_0_w22;  // <1,0>
  float_24_8                    biasIn_0_w23;  // <1,0>
  float_24_8                    biasIn_0_w24;  // <1,0>
  float_24_8                    biasIn_0_w25;  // <1,0>
  float_24_8                    biasIn_0_w26;  // <1,0>
  float_24_8                    biasIn_0_w27;  // <1,0>
  float_24_8                    biasIn_0_w28;  // <1,0>
  float_24_8                    biasIn_0_w29;  // <1,0>
  float_24_8                    biasIn_0_w3;  // <1,0>
  float_24_8                    biasIn_0_w30;  // <1,0>
  float_24_8                    biasIn_0_w31;  // <1,0>
  float_24_8                    biasIn_0_w32;  // <1,0>
  float_24_8                    biasIn_0_w33;  // <1,0>
  float_24_8                    biasIn_0_w34;  // <1,0>
  float_24_8                    biasIn_0_w35;  // <1,0>
  float_24_8                    biasIn_0_w36;  // <1,0>
  float_24_8                    biasIn_0_w37;  // <1,0>
  float_24_8                    biasIn_0_w38;  // <1,0>
  float_24_8                    biasIn_0_w39;  // <1,0>
  float_24_8                    biasIn_0_w4;  // <1,0>
  float_24_8                    biasIn_0_w40;  // <1,0>
  float_24_8                    biasIn_0_w41;  // <1,0>
  float_24_8                    biasIn_0_w42;  // <1,0>
  float_24_8                    biasIn_0_w43;  // <1,0>
  float_24_8                    biasIn_0_w44;  // <1,0>
  float_24_8                    biasIn_0_w45;  // <1,0>
  float_24_8                    biasIn_0_w46;  // <1,0>
  float_24_8                    biasIn_0_w47;  // <1,0>
  float_24_8                    biasIn_0_w48;  // <1,0>
  float_24_8                    biasIn_0_w49;  // <1,0>
  float_24_8                    biasIn_0_w5;  // <1,0>
  float_24_8                    biasIn_0_w50;  // <1,0>
  float_24_8                    biasIn_0_w51;  // <1,0>
  float_24_8                    biasIn_0_w52;  // <1,0>
  float_24_8                    biasIn_0_w53;  // <1,0>
  float_24_8                    biasIn_0_w54;  // <1,0>
  float_24_8                    biasIn_0_w55;  // <1,0>
  float_24_8                    biasIn_0_w56;  // <1,0>
  float_24_8                    biasIn_0_w57;  // <1,0>
  float_24_8                    biasIn_0_w58;  // <1,0>
  float_24_8                    biasIn_0_w59;  // <1,0>
  float_24_8                    biasIn_0_w6;  // <1,0>
  float_24_8                    biasIn_0_w60;  // <1,0>
  float_24_8                    biasIn_0_w61;  // <1,0>
  float_24_8                    biasIn_0_w62;  // <1,0>
  float_24_8                    biasIn_0_w63;  // <1,0>
  float_24_8                    biasIn_0_w64;  // <1,0>
  float_24_8                    biasIn_0_w65;  // <1,0>
  float_24_8                    biasIn_0_w66;  // <1,0>
  float_24_8                    biasIn_0_w67;  // <1,0>
  float_24_8                    biasIn_0_w68;  // <1,0>
  float_24_8                    biasIn_0_w69;  // <1,0>
  float_24_8                    biasIn_0_w7;  // <1,0>
  float_24_8                    biasIn_0_w70;  // <1,0>
  float_24_8                    biasIn_0_w71;  // <1,0>
  float_24_8                    biasIn_0_w72;  // <1,0>
  float_24_8                    biasIn_0_w73;  // <1,0>
  float_24_8                    biasIn_0_w74;  // <1,0>
  float_24_8                    biasIn_0_w75;  // <1,0>
  float_24_8                    biasIn_0_w76;  // <1,0>
  float_24_8                    biasIn_0_w77;  // <1,0>
  float_24_8                    biasIn_0_w78;  // <1,0>
  float_24_8                    biasIn_0_w79;  // <1,0>
  float_24_8                    biasIn_0_w8;  // <1,0>
  float_24_8                    biasIn_0_w80;  // <1,0>
  float_24_8                    biasIn_0_w81;  // <1,0>
  float_24_8                    biasIn_0_w82;  // <1,0>
  float_24_8                    biasIn_0_w83;  // <1,0>
  float_24_8                    biasIn_0_w84;  // <1,0>
  float_24_8                    biasIn_0_w85;  // <1,0>
  float_24_8                    biasIn_0_w86;  // <1,0>
  float_24_8                    biasIn_0_w87;  // <1,0>
  float_24_8                    biasIn_0_w88;  // <1,0>
  float_24_8                    biasIn_0_w89;  // <1,0>
  float_24_8                    biasIn_0_w9;  // <1,0>
  float_24_8                    biasIn_0_w90;  // <1,0>
  float_24_8                    biasIn_0_w91;  // <1,0>
  float_24_8                    biasIn_0_w92;  // <1,0>
  float_24_8                    biasIn_0_w93;  // <1,0>
  float_24_8                    biasIn_0_w94;  // <1,0>
  float_24_8                    biasIn_0_w95;  // <1,0>
  float_24_8                    biasIn_0_w96;  // <1,0>
  float_24_8                    biasIn_0_w97;  // <1,0>
  float_24_8                    biasIn_0_w98;  // <1,0>
  float_24_8                    biasIn_0_w99;  // <1,0>
  float_24_8                    wireOut_w0;  // <1,0>
  float_24_8                    wireOut_w1;  // <1,0>
  float_24_8                    wireOut_w10;  // <1,0>
  float_24_8                    wireOut_w100;  // <1,0>
  float_24_8                    wireOut_w101;  // <1,0>
  float_24_8                    wireOut_w102;  // <1,0>
  float_24_8                    wireOut_w103;  // <1,0>
  float_24_8                    wireOut_w104;  // <1,0>
  float_24_8                    wireOut_w105;  // <1,0>
  float_24_8                    wireOut_w106;  // <1,0>
  float_24_8                    wireOut_w107;  // <1,0>
  float_24_8                    wireOut_w108;  // <1,0>
  float_24_8                    wireOut_w109;  // <1,0>
  float_24_8                    wireOut_w11;  // <1,0>
  float_24_8                    wireOut_w110;  // <1,0>
  float_24_8                    wireOut_w111;  // <1,0>
  float_24_8                    wireOut_w112;  // <1,0>
  float_24_8                    wireOut_w113;  // <1,0>
  float_24_8                    wireOut_w114;  // <1,0>
  float_24_8                    wireOut_w115;  // <1,0>
  float_24_8                    wireOut_w116;  // <1,0>
  float_24_8                    wireOut_w117;  // <1,0>
  float_24_8                    wireOut_w118;  // <1,0>
  float_24_8                    wireOut_w119;  // <1,0>
  float_24_8                    wireOut_w12;  // <1,0>
  float_24_8                    wireOut_w120;  // <1,0>
  float_24_8                    wireOut_w121;  // <1,0>
  float_24_8                    wireOut_w122;  // <1,0>
  float_24_8                    wireOut_w123;  // <1,0>
  float_24_8                    wireOut_w124;  // <1,0>
  float_24_8                    wireOut_w125;  // <1,0>
  float_24_8                    wireOut_w126;  // <1,0>
  float_24_8                    wireOut_w127;  // <1,0>
  float_24_8                    wireOut_w13;  // <1,0>
  float_24_8                    wireOut_w14;  // <1,0>
  float_24_8                    wireOut_w15;  // <1,0>
  float_24_8                    wireOut_w16;  // <1,0>
  float_24_8                    wireOut_w17;  // <1,0>
  float_24_8                    wireOut_w18;  // <1,0>
  float_24_8                    wireOut_w19;  // <1,0>
  float_24_8                    wireOut_w2;  // <1,0>
  float_24_8                    wireOut_w20;  // <1,0>
  float_24_8                    wireOut_w21;  // <1,0>
  float_24_8                    wireOut_w22;  // <1,0>
  float_24_8                    wireOut_w23;  // <1,0>
  float_24_8                    wireOut_w24;  // <1,0>
  float_24_8                    wireOut_w25;  // <1,0>
  float_24_8                    wireOut_w26;  // <1,0>
  float_24_8                    wireOut_w27;  // <1,0>
  float_24_8                    wireOut_w28;  // <1,0>
  float_24_8                    wireOut_w29;  // <1,0>
  float_24_8                    wireOut_w3;  // <1,0>
  float_24_8                    wireOut_w30;  // <1,0>
  float_24_8                    wireOut_w31;  // <1,0>
  float_24_8                    wireOut_w32;  // <1,0>
  float_24_8                    wireOut_w33;  // <1,0>
  float_24_8                    wireOut_w34;  // <1,0>
  float_24_8                    wireOut_w35;  // <1,0>
  float_24_8                    wireOut_w36;  // <1,0>
  float_24_8                    wireOut_w37;  // <1,0>
  float_24_8                    wireOut_w38;  // <1,0>
  float_24_8                    wireOut_w39;  // <1,0>
  float_24_8                    wireOut_w4;  // <1,0>
  float_24_8                    wireOut_w40;  // <1,0>
  float_24_8                    wireOut_w41;  // <1,0>
  float_24_8                    wireOut_w42;  // <1,0>
  float_24_8                    wireOut_w43;  // <1,0>
  float_24_8                    wireOut_w44;  // <1,0>
  float_24_8                    wireOut_w45;  // <1,0>
  float_24_8                    wireOut_w46;  // <1,0>
  float_24_8                    wireOut_w47;  // <1,0>
  float_24_8                    wireOut_w48;  // <1,0>
  float_24_8                    wireOut_w49;  // <1,0>
  float_24_8                    wireOut_w5;  // <1,0>
  float_24_8                    wireOut_w50;  // <1,0>
  float_24_8                    wireOut_w51;  // <1,0>
  float_24_8                    wireOut_w52;  // <1,0>
  float_24_8                    wireOut_w53;  // <1,0>
  float_24_8                    wireOut_w54;  // <1,0>
  float_24_8                    wireOut_w55;  // <1,0>
  float_24_8                    wireOut_w56;  // <1,0>
  float_24_8                    wireOut_w57;  // <1,0>
  float_24_8                    wireOut_w58;  // <1,0>
  float_24_8                    wireOut_w59;  // <1,0>
  float_24_8                    wireOut_w6;  // <1,0>
  float_24_8                    wireOut_w60;  // <1,0>
  float_24_8                    wireOut_w61;  // <1,0>
  float_24_8                    wireOut_w62;  // <1,0>
  float_24_8                    wireOut_w63;  // <1,0>
  float_24_8                    wireOut_w64;  // <1,0>
  float_24_8                    wireOut_w65;  // <1,0>
  float_24_8                    wireOut_w66;  // <1,0>
  float_24_8                    wireOut_w67;  // <1,0>
  float_24_8                    wireOut_w68;  // <1,0>
  float_24_8                    wireOut_w69;  // <1,0>
  float_24_8                    wireOut_w7;  // <1,0>
  float_24_8                    wireOut_w70;  // <1,0>
  float_24_8                    wireOut_w71;  // <1,0>
  float_24_8                    wireOut_w72;  // <1,0>
  float_24_8                    wireOut_w73;  // <1,0>
  float_24_8                    wireOut_w74;  // <1,0>
  float_24_8                    wireOut_w75;  // <1,0>
  float_24_8                    wireOut_w76;  // <1,0>
  float_24_8                    wireOut_w77;  // <1,0>
  float_24_8                    wireOut_w78;  // <1,0>
  float_24_8                    wireOut_w79;  // <1,0>
  float_24_8                    wireOut_w8;  // <1,0>
  float_24_8                    wireOut_w80;  // <1,0>
  float_24_8                    wireOut_w81;  // <1,0>
  float_24_8                    wireOut_w82;  // <1,0>
  float_24_8                    wireOut_w83;  // <1,0>
  float_24_8                    wireOut_w84;  // <1,0>
  float_24_8                    wireOut_w85;  // <1,0>
  float_24_8                    wireOut_w86;  // <1,0>
  float_24_8                    wireOut_w87;  // <1,0>
  float_24_8                    wireOut_w88;  // <1,0>
  float_24_8                    wireOut_w89;  // <1,0>
  float_24_8                    wireOut_w9;  // <1,0>
  float_24_8                    wireOut_w90;  // <1,0>
  float_24_8                    wireOut_w91;  // <1,0>
  float_24_8                    wireOut_w92;  // <1,0>
  float_24_8                    wireOut_w93;  // <1,0>
  float_24_8                    wireOut_w94;  // <1,0>
  float_24_8                    wireOut_w95;  // <1,0>
  float_24_8                    wireOut_w96;  // <1,0>
  float_24_8                    wireOut_w97;  // <1,0>
  float_24_8                    wireOut_w98;  // <1,0>
  float_24_8                    wireOut_w99;  // <1,0>


// Registers 

  float_24_8                    biasIn_0_r1;  // <1,0>
  float_24_8                    biasIn_0_r10;  // <1,0>
  float_24_8                    biasIn_0_r100;  // <1,0>
  float_24_8                    biasIn_0_r101;  // <1,0>
  float_24_8                    biasIn_0_r102;  // <1,0>
  float_24_8                    biasIn_0_r103;  // <1,0>
  float_24_8                    biasIn_0_r104;  // <1,0>
  float_24_8                    biasIn_0_r105;  // <1,0>
  float_24_8                    biasIn_0_r106;  // <1,0>
  float_24_8                    biasIn_0_r107;  // <1,0>
  float_24_8                    biasIn_0_r108;  // <1,0>
  float_24_8                    biasIn_0_r109;  // <1,0>
  float_24_8                    biasIn_0_r11;  // <1,0>
  float_24_8                    biasIn_0_r110;  // <1,0>
  float_24_8                    biasIn_0_r111;  // <1,0>
  float_24_8                    biasIn_0_r112;  // <1,0>
  float_24_8                    biasIn_0_r113;  // <1,0>
  float_24_8                    biasIn_0_r114;  // <1,0>
  float_24_8                    biasIn_0_r115;  // <1,0>
  float_24_8                    biasIn_0_r116;  // <1,0>
  float_24_8                    biasIn_0_r117;  // <1,0>
  float_24_8                    biasIn_0_r118;  // <1,0>
  float_24_8                    biasIn_0_r119;  // <1,0>
  float_24_8                    biasIn_0_r12;  // <1,0>
  float_24_8                    biasIn_0_r120;  // <1,0>
  float_24_8                    biasIn_0_r121;  // <1,0>
  float_24_8                    biasIn_0_r122;  // <1,0>
  float_24_8                    biasIn_0_r123;  // <1,0>
  float_24_8                    biasIn_0_r124;  // <1,0>
  float_24_8                    biasIn_0_r125;  // <1,0>
  float_24_8                    biasIn_0_r126;  // <1,0>
  float_24_8                    biasIn_0_r127;  // <1,0>
  float_24_8                    biasIn_0_r128;  // <1,0>
  float_24_8                    biasIn_0_r13;  // <1,0>
  float_24_8                    biasIn_0_r14;  // <1,0>
  float_24_8                    biasIn_0_r15;  // <1,0>
  float_24_8                    biasIn_0_r16;  // <1,0>
  float_24_8                    biasIn_0_r17;  // <1,0>
  float_24_8                    biasIn_0_r18;  // <1,0>
  float_24_8                    biasIn_0_r19;  // <1,0>
  float_24_8                    biasIn_0_r2;  // <1,0>
  float_24_8                    biasIn_0_r20;  // <1,0>
  float_24_8                    biasIn_0_r21;  // <1,0>
  float_24_8                    biasIn_0_r22;  // <1,0>
  float_24_8                    biasIn_0_r23;  // <1,0>
  float_24_8                    biasIn_0_r24;  // <1,0>
  float_24_8                    biasIn_0_r25;  // <1,0>
  float_24_8                    biasIn_0_r26;  // <1,0>
  float_24_8                    biasIn_0_r27;  // <1,0>
  float_24_8                    biasIn_0_r28;  // <1,0>
  float_24_8                    biasIn_0_r29;  // <1,0>
  float_24_8                    biasIn_0_r3;  // <1,0>
  float_24_8                    biasIn_0_r30;  // <1,0>
  float_24_8                    biasIn_0_r31;  // <1,0>
  float_24_8                    biasIn_0_r32;  // <1,0>
  float_24_8                    biasIn_0_r33;  // <1,0>
  float_24_8                    biasIn_0_r34;  // <1,0>
  float_24_8                    biasIn_0_r35;  // <1,0>
  float_24_8                    biasIn_0_r36;  // <1,0>
  float_24_8                    biasIn_0_r37;  // <1,0>
  float_24_8                    biasIn_0_r38;  // <1,0>
  float_24_8                    biasIn_0_r39;  // <1,0>
  float_24_8                    biasIn_0_r4;  // <1,0>
  float_24_8                    biasIn_0_r40;  // <1,0>
  float_24_8                    biasIn_0_r41;  // <1,0>
  float_24_8                    biasIn_0_r42;  // <1,0>
  float_24_8                    biasIn_0_r43;  // <1,0>
  float_24_8                    biasIn_0_r44;  // <1,0>
  float_24_8                    biasIn_0_r45;  // <1,0>
  float_24_8                    biasIn_0_r46;  // <1,0>
  float_24_8                    biasIn_0_r47;  // <1,0>
  float_24_8                    biasIn_0_r48;  // <1,0>
  float_24_8                    biasIn_0_r49;  // <1,0>
  float_24_8                    biasIn_0_r5;  // <1,0>
  float_24_8                    biasIn_0_r50;  // <1,0>
  float_24_8                    biasIn_0_r51;  // <1,0>
  float_24_8                    biasIn_0_r52;  // <1,0>
  float_24_8                    biasIn_0_r53;  // <1,0>
  float_24_8                    biasIn_0_r54;  // <1,0>
  float_24_8                    biasIn_0_r55;  // <1,0>
  float_24_8                    biasIn_0_r56;  // <1,0>
  float_24_8                    biasIn_0_r57;  // <1,0>
  float_24_8                    biasIn_0_r58;  // <1,0>
  float_24_8                    biasIn_0_r59;  // <1,0>
  float_24_8                    biasIn_0_r6;  // <1,0>
  float_24_8                    biasIn_0_r60;  // <1,0>
  float_24_8                    biasIn_0_r61;  // <1,0>
  float_24_8                    biasIn_0_r62;  // <1,0>
  float_24_8                    biasIn_0_r63;  // <1,0>
  float_24_8                    biasIn_0_r64;  // <1,0>
  float_24_8                    biasIn_0_r65;  // <1,0>
  float_24_8                    biasIn_0_r66;  // <1,0>
  float_24_8                    biasIn_0_r67;  // <1,0>
  float_24_8                    biasIn_0_r68;  // <1,0>
  float_24_8                    biasIn_0_r69;  // <1,0>
  float_24_8                    biasIn_0_r7;  // <1,0>
  float_24_8                    biasIn_0_r70;  // <1,0>
  float_24_8                    biasIn_0_r71;  // <1,0>
  float_24_8                    biasIn_0_r72;  // <1,0>
  float_24_8                    biasIn_0_r73;  // <1,0>
  float_24_8                    biasIn_0_r74;  // <1,0>
  float_24_8                    biasIn_0_r75;  // <1,0>
  float_24_8                    biasIn_0_r76;  // <1,0>
  float_24_8                    biasIn_0_r77;  // <1,0>
  float_24_8                    biasIn_0_r78;  // <1,0>
  float_24_8                    biasIn_0_r79;  // <1,0>
  float_24_8                    biasIn_0_r8;  // <1,0>
  float_24_8                    biasIn_0_r80;  // <1,0>
  float_24_8                    biasIn_0_r81;  // <1,0>
  float_24_8                    biasIn_0_r82;  // <1,0>
  float_24_8                    biasIn_0_r83;  // <1,0>
  float_24_8                    biasIn_0_r84;  // <1,0>
  float_24_8                    biasIn_0_r85;  // <1,0>
  float_24_8                    biasIn_0_r86;  // <1,0>
  float_24_8                    biasIn_0_r87;  // <1,0>
  float_24_8                    biasIn_0_r88;  // <1,0>
  float_24_8                    biasIn_0_r89;  // <1,0>
  float_24_8                    biasIn_0_r9;  // <1,0>
  float_24_8                    biasIn_0_r90;  // <1,0>
  float_24_8                    biasIn_0_r91;  // <1,0>
  float_24_8                    biasIn_0_r92;  // <1,0>
  float_24_8                    biasIn_0_r93;  // <1,0>
  float_24_8                    biasIn_0_r94;  // <1,0>
  float_24_8                    biasIn_0_r95;  // <1,0>
  float_24_8                    biasIn_0_r96;  // <1,0>
  float_24_8                    biasIn_0_r97;  // <1,0>
  float_24_8                    biasIn_0_r98;  // <1,0>
  float_24_8                    biasIn_0_r99;  // <1,0>
  float_24_8                    outLine_w0;  // <1,0>
  float_24_8                    outLine_w1;  // <1,0>
  float_24_8                    outLine_w10;  // <1,0>
  float_24_8                    outLine_w100;  // <1,0>
  float_24_8                    outLine_w101;  // <1,0>
  float_24_8                    outLine_w102;  // <1,0>
  float_24_8                    outLine_w103;  // <1,0>
  float_24_8                    outLine_w104;  // <1,0>
  float_24_8                    outLine_w105;  // <1,0>
  float_24_8                    outLine_w106;  // <1,0>
  float_24_8                    outLine_w107;  // <1,0>
  float_24_8                    outLine_w108;  // <1,0>
  float_24_8                    outLine_w109;  // <1,0>
  float_24_8                    outLine_w11;  // <1,0>
  float_24_8                    outLine_w110;  // <1,0>
  float_24_8                    outLine_w111;  // <1,0>
  float_24_8                    outLine_w112;  // <1,0>
  float_24_8                    outLine_w113;  // <1,0>
  float_24_8                    outLine_w114;  // <1,0>
  float_24_8                    outLine_w115;  // <1,0>
  float_24_8                    outLine_w116;  // <1,0>
  float_24_8                    outLine_w117;  // <1,0>
  float_24_8                    outLine_w118;  // <1,0>
  float_24_8                    outLine_w119;  // <1,0>
  float_24_8                    outLine_w12;  // <1,0>
  float_24_8                    outLine_w120;  // <1,0>
  float_24_8                    outLine_w121;  // <1,0>
  float_24_8                    outLine_w122;  // <1,0>
  float_24_8                    outLine_w123;  // <1,0>
  float_24_8                    outLine_w124;  // <1,0>
  float_24_8                    outLine_w125;  // <1,0>
  float_24_8                    outLine_w126;  // <1,0>
  float_24_8                    outLine_w127;  // <1,0>
  float_24_8                    outLine_w13;  // <1,0>
  float_24_8                    outLine_w14;  // <1,0>
  float_24_8                    outLine_w15;  // <1,0>
  float_24_8                    outLine_w16;  // <1,0>
  float_24_8                    outLine_w17;  // <1,0>
  float_24_8                    outLine_w18;  // <1,0>
  float_24_8                    outLine_w19;  // <1,0>
  float_24_8                    outLine_w2;  // <1,0>
  float_24_8                    outLine_w20;  // <1,0>
  float_24_8                    outLine_w21;  // <1,0>
  float_24_8                    outLine_w22;  // <1,0>
  float_24_8                    outLine_w23;  // <1,0>
  float_24_8                    outLine_w24;  // <1,0>
  float_24_8                    outLine_w25;  // <1,0>
  float_24_8                    outLine_w26;  // <1,0>
  float_24_8                    outLine_w27;  // <1,0>
  float_24_8                    outLine_w28;  // <1,0>
  float_24_8                    outLine_w29;  // <1,0>
  float_24_8                    outLine_w3;  // <1,0>
  float_24_8                    outLine_w30;  // <1,0>
  float_24_8                    outLine_w31;  // <1,0>
  float_24_8                    outLine_w32;  // <1,0>
  float_24_8                    outLine_w33;  // <1,0>
  float_24_8                    outLine_w34;  // <1,0>
  float_24_8                    outLine_w35;  // <1,0>
  float_24_8                    outLine_w36;  // <1,0>
  float_24_8                    outLine_w37;  // <1,0>
  float_24_8                    outLine_w38;  // <1,0>
  float_24_8                    outLine_w39;  // <1,0>
  float_24_8                    outLine_w4;  // <1,0>
  float_24_8                    outLine_w40;  // <1,0>
  float_24_8                    outLine_w41;  // <1,0>
  float_24_8                    outLine_w42;  // <1,0>
  float_24_8                    outLine_w43;  // <1,0>
  float_24_8                    outLine_w44;  // <1,0>
  float_24_8                    outLine_w45;  // <1,0>
  float_24_8                    outLine_w46;  // <1,0>
  float_24_8                    outLine_w47;  // <1,0>
  float_24_8                    outLine_w48;  // <1,0>
  float_24_8                    outLine_w49;  // <1,0>
  float_24_8                    outLine_w5;  // <1,0>
  float_24_8                    outLine_w50;  // <1,0>
  float_24_8                    outLine_w51;  // <1,0>
  float_24_8                    outLine_w52;  // <1,0>
  float_24_8                    outLine_w53;  // <1,0>
  float_24_8                    outLine_w54;  // <1,0>
  float_24_8                    outLine_w55;  // <1,0>
  float_24_8                    outLine_w56;  // <1,0>
  float_24_8                    outLine_w57;  // <1,0>
  float_24_8                    outLine_w58;  // <1,0>
  float_24_8                    outLine_w59;  // <1,0>
  float_24_8                    outLine_w6;  // <1,0>
  float_24_8                    outLine_w60;  // <1,0>
  float_24_8                    outLine_w61;  // <1,0>
  float_24_8                    outLine_w62;  // <1,0>
  float_24_8                    outLine_w63;  // <1,0>
  float_24_8                    outLine_w64;  // <1,0>
  float_24_8                    outLine_w65;  // <1,0>
  float_24_8                    outLine_w66;  // <1,0>
  float_24_8                    outLine_w67;  // <1,0>
  float_24_8                    outLine_w68;  // <1,0>
  float_24_8                    outLine_w69;  // <1,0>
  float_24_8                    outLine_w7;  // <1,0>
  float_24_8                    outLine_w70;  // <1,0>
  float_24_8                    outLine_w71;  // <1,0>
  float_24_8                    outLine_w72;  // <1,0>
  float_24_8                    outLine_w73;  // <1,0>
  float_24_8                    outLine_w74;  // <1,0>
  float_24_8                    outLine_w75;  // <1,0>
  float_24_8                    outLine_w76;  // <1,0>
  float_24_8                    outLine_w77;  // <1,0>
  float_24_8                    outLine_w78;  // <1,0>
  float_24_8                    outLine_w79;  // <1,0>
  float_24_8                    outLine_w8;  // <1,0>
  float_24_8                    outLine_w80;  // <1,0>
  float_24_8                    outLine_w81;  // <1,0>
  float_24_8                    outLine_w82;  // <1,0>
  float_24_8                    outLine_w83;  // <1,0>
  float_24_8                    outLine_w84;  // <1,0>
  float_24_8                    outLine_w85;  // <1,0>
  float_24_8                    outLine_w86;  // <1,0>
  float_24_8                    outLine_w87;  // <1,0>
  float_24_8                    outLine_w88;  // <1,0>
  float_24_8                    outLine_w89;  // <1,0>
  float_24_8                    outLine_w9;  // <1,0>
  float_24_8                    outLine_w90;  // <1,0>
  float_24_8                    outLine_w91;  // <1,0>
  float_24_8                    outLine_w92;  // <1,0>
  float_24_8                    outLine_w93;  // <1,0>
  float_24_8                    outLine_w94;  // <1,0>
  float_24_8                    outLine_w95;  // <1,0>
  float_24_8                    outLine_w96;  // <1,0>
  float_24_8                    outLine_w97;  // <1,0>
  float_24_8                    outLine_w98;  // <1,0>
  float_24_8                    outLine_w99;  // <1,0>
  reg                           valid0            ;  // <1,0>
  reg                           valid1            ;  // <1,0>


// Other



always @(posedge clk) begin
  if (reset) begin
    biasIn_0_r1 <= 'd0;
    biasIn_0_r2 <= 'd0;
    biasIn_0_r3 <= 'd0;
    biasIn_0_r4 <= 'd0;
    biasIn_0_r5 <= 'd0;
    biasIn_0_r6 <= 'd0;
    biasIn_0_r7 <= 'd0;
    biasIn_0_r8 <= 'd0;
    biasIn_0_r9 <= 'd0;
    biasIn_0_r10 <= 'd0;
    biasIn_0_r11 <= 'd0;
    biasIn_0_r12 <= 'd0;
    biasIn_0_r13 <= 'd0;
    biasIn_0_r14 <= 'd0;
    biasIn_0_r15 <= 'd0;
    biasIn_0_r16 <= 'd0;
    biasIn_0_r17 <= 'd0;
    biasIn_0_r18 <= 'd0;
    biasIn_0_r19 <= 'd0;
    biasIn_0_r20 <= 'd0;
    biasIn_0_r21 <= 'd0;
    biasIn_0_r22 <= 'd0;
    biasIn_0_r23 <= 'd0;
    biasIn_0_r24 <= 'd0;
    biasIn_0_r25 <= 'd0;
    biasIn_0_r26 <= 'd0;
    biasIn_0_r27 <= 'd0;
    biasIn_0_r28 <= 'd0;
    biasIn_0_r29 <= 'd0;
    biasIn_0_r30 <= 'd0;
    biasIn_0_r31 <= 'd0;
    biasIn_0_r32 <= 'd0;
    biasIn_0_r33 <= 'd0;
    biasIn_0_r34 <= 'd0;
    biasIn_0_r35 <= 'd0;
    biasIn_0_r36 <= 'd0;
    biasIn_0_r37 <= 'd0;
    biasIn_0_r38 <= 'd0;
    biasIn_0_r39 <= 'd0;
    biasIn_0_r40 <= 'd0;
    biasIn_0_r41 <= 'd0;
    biasIn_0_r42 <= 'd0;
    biasIn_0_r43 <= 'd0;
    biasIn_0_r44 <= 'd0;
    biasIn_0_r45 <= 'd0;
    biasIn_0_r46 <= 'd0;
    biasIn_0_r47 <= 'd0;
    biasIn_0_r48 <= 'd0;
    biasIn_0_r49 <= 'd0;
    biasIn_0_r50 <= 'd0;
    biasIn_0_r51 <= 'd0;
    biasIn_0_r52 <= 'd0;
    biasIn_0_r53 <= 'd0;
    biasIn_0_r54 <= 'd0;
    biasIn_0_r55 <= 'd0;
    biasIn_0_r56 <= 'd0;
    biasIn_0_r57 <= 'd0;
    biasIn_0_r58 <= 'd0;
    biasIn_0_r59 <= 'd0;
    biasIn_0_r60 <= 'd0;
    biasIn_0_r61 <= 'd0;
    biasIn_0_r62 <= 'd0;
    biasIn_0_r63 <= 'd0;
    biasIn_0_r64 <= 'd0;
    biasIn_0_r65 <= 'd0;
    biasIn_0_r66 <= 'd0;
    biasIn_0_r67 <= 'd0;
    biasIn_0_r68 <= 'd0;
    biasIn_0_r69 <= 'd0;
    biasIn_0_r70 <= 'd0;
    biasIn_0_r71 <= 'd0;
    biasIn_0_r72 <= 'd0;
    biasIn_0_r73 <= 'd0;
    biasIn_0_r74 <= 'd0;
    biasIn_0_r75 <= 'd0;
    biasIn_0_r76 <= 'd0;
    biasIn_0_r77 <= 'd0;
    biasIn_0_r78 <= 'd0;
    biasIn_0_r79 <= 'd0;
    biasIn_0_r80 <= 'd0;
    biasIn_0_r81 <= 'd0;
    biasIn_0_r82 <= 'd0;
    biasIn_0_r83 <= 'd0;
    biasIn_0_r84 <= 'd0;
    biasIn_0_r85 <= 'd0;
    biasIn_0_r86 <= 'd0;
    biasIn_0_r87 <= 'd0;
    biasIn_0_r88 <= 'd0;
    biasIn_0_r89 <= 'd0;
    biasIn_0_r90 <= 'd0;
    biasIn_0_r91 <= 'd0;
    biasIn_0_r92 <= 'd0;
    biasIn_0_r93 <= 'd0;
    biasIn_0_r94 <= 'd0;
    biasIn_0_r95 <= 'd0;
    biasIn_0_r96 <= 'd0;
    biasIn_0_r97 <= 'd0;
    biasIn_0_r98 <= 'd0;
    biasIn_0_r99 <= 'd0;
    biasIn_0_r100 <= 'd0;
    biasIn_0_r101 <= 'd0;
    biasIn_0_r102 <= 'd0;
    biasIn_0_r103 <= 'd0;
    biasIn_0_r104 <= 'd0;
    biasIn_0_r105 <= 'd0;
    biasIn_0_r106 <= 'd0;
    biasIn_0_r107 <= 'd0;
    biasIn_0_r108 <= 'd0;
    biasIn_0_r109 <= 'd0;
    biasIn_0_r110 <= 'd0;
    biasIn_0_r111 <= 'd0;
    biasIn_0_r112 <= 'd0;
    biasIn_0_r113 <= 'd0;
    biasIn_0_r114 <= 'd0;
    biasIn_0_r115 <= 'd0;
    biasIn_0_r116 <= 'd0;
    biasIn_0_r117 <= 'd0;
    biasIn_0_r118 <= 'd0;
    biasIn_0_r119 <= 'd0;
    biasIn_0_r120 <= 'd0;
    biasIn_0_r121 <= 'd0;
    biasIn_0_r122 <= 'd0;
    biasIn_0_r123 <= 'd0;
    biasIn_0_r124 <= 'd0;
    biasIn_0_r125 <= 'd0;
    biasIn_0_r126 <= 'd0;
    biasIn_0_r127 <= 'd0;
    biasIn_0_r128 <= 'd0;
  end
  else begin
    biasIn_0_r1 <= biasIn_0;
    biasIn_0_r2 <= biasIn_0_r1;
    biasIn_0_r3 <= biasIn_0_r2;
    biasIn_0_r4 <= biasIn_0_r3;
    biasIn_0_r5 <= biasIn_0_r4;
    biasIn_0_r6 <= biasIn_0_r5;
    biasIn_0_r7 <= biasIn_0_r6;
    biasIn_0_r8 <= biasIn_0_r7;
    biasIn_0_r9 <= biasIn_0_r8;
    biasIn_0_r10 <= biasIn_0_r9;
    biasIn_0_r11 <= biasIn_0_r10;
    biasIn_0_r12 <= biasIn_0_r11;
    biasIn_0_r13 <= biasIn_0_r12;
    biasIn_0_r14 <= biasIn_0_r13;
    biasIn_0_r15 <= biasIn_0_r14;
    biasIn_0_r16 <= biasIn_0_r15;
    biasIn_0_r17 <= biasIn_0_r16;
    biasIn_0_r18 <= biasIn_0_r17;
    biasIn_0_r19 <= biasIn_0_r18;
    biasIn_0_r20 <= biasIn_0_r19;
    biasIn_0_r21 <= biasIn_0_r20;
    biasIn_0_r22 <= biasIn_0_r21;
    biasIn_0_r23 <= biasIn_0_r22;
    biasIn_0_r24 <= biasIn_0_r23;
    biasIn_0_r25 <= biasIn_0_r24;
    biasIn_0_r26 <= biasIn_0_r25;
    biasIn_0_r27 <= biasIn_0_r26;
    biasIn_0_r28 <= biasIn_0_r27;
    biasIn_0_r29 <= biasIn_0_r28;
    biasIn_0_r30 <= biasIn_0_r29;
    biasIn_0_r31 <= biasIn_0_r30;
    biasIn_0_r32 <= biasIn_0_r31;
    biasIn_0_r33 <= biasIn_0_r32;
    biasIn_0_r34 <= biasIn_0_r33;
    biasIn_0_r35 <= biasIn_0_r34;
    biasIn_0_r36 <= biasIn_0_r35;
    biasIn_0_r37 <= biasIn_0_r36;
    biasIn_0_r38 <= biasIn_0_r37;
    biasIn_0_r39 <= biasIn_0_r38;
    biasIn_0_r40 <= biasIn_0_r39;
    biasIn_0_r41 <= biasIn_0_r40;
    biasIn_0_r42 <= biasIn_0_r41;
    biasIn_0_r43 <= biasIn_0_r42;
    biasIn_0_r44 <= biasIn_0_r43;
    biasIn_0_r45 <= biasIn_0_r44;
    biasIn_0_r46 <= biasIn_0_r45;
    biasIn_0_r47 <= biasIn_0_r46;
    biasIn_0_r48 <= biasIn_0_r47;
    biasIn_0_r49 <= biasIn_0_r48;
    biasIn_0_r50 <= biasIn_0_r49;
    biasIn_0_r51 <= biasIn_0_r50;
    biasIn_0_r52 <= biasIn_0_r51;
    biasIn_0_r53 <= biasIn_0_r52;
    biasIn_0_r54 <= biasIn_0_r53;
    biasIn_0_r55 <= biasIn_0_r54;
    biasIn_0_r56 <= biasIn_0_r55;
    biasIn_0_r57 <= biasIn_0_r56;
    biasIn_0_r58 <= biasIn_0_r57;
    biasIn_0_r59 <= biasIn_0_r58;
    biasIn_0_r60 <= biasIn_0_r59;
    biasIn_0_r61 <= biasIn_0_r60;
    biasIn_0_r62 <= biasIn_0_r61;
    biasIn_0_r63 <= biasIn_0_r62;
    biasIn_0_r64 <= biasIn_0_r63;
    biasIn_0_r65 <= biasIn_0_r64;
    biasIn_0_r66 <= biasIn_0_r65;
    biasIn_0_r67 <= biasIn_0_r66;
    biasIn_0_r68 <= biasIn_0_r67;
    biasIn_0_r69 <= biasIn_0_r68;
    biasIn_0_r70 <= biasIn_0_r69;
    biasIn_0_r71 <= biasIn_0_r70;
    biasIn_0_r72 <= biasIn_0_r71;
    biasIn_0_r73 <= biasIn_0_r72;
    biasIn_0_r74 <= biasIn_0_r73;
    biasIn_0_r75 <= biasIn_0_r74;
    biasIn_0_r76 <= biasIn_0_r75;
    biasIn_0_r77 <= biasIn_0_r76;
    biasIn_0_r78 <= biasIn_0_r77;
    biasIn_0_r79 <= biasIn_0_r78;
    biasIn_0_r80 <= biasIn_0_r79;
    biasIn_0_r81 <= biasIn_0_r80;
    biasIn_0_r82 <= biasIn_0_r81;
    biasIn_0_r83 <= biasIn_0_r82;
    biasIn_0_r84 <= biasIn_0_r83;
    biasIn_0_r85 <= biasIn_0_r84;
    biasIn_0_r86 <= biasIn_0_r85;
    biasIn_0_r87 <= biasIn_0_r86;
    biasIn_0_r88 <= biasIn_0_r87;
    biasIn_0_r89 <= biasIn_0_r88;
    biasIn_0_r90 <= biasIn_0_r89;
    biasIn_0_r91 <= biasIn_0_r90;
    biasIn_0_r92 <= biasIn_0_r91;
    biasIn_0_r93 <= biasIn_0_r92;
    biasIn_0_r94 <= biasIn_0_r93;
    biasIn_0_r95 <= biasIn_0_r94;
    biasIn_0_r96 <= biasIn_0_r95;
    biasIn_0_r97 <= biasIn_0_r96;
    biasIn_0_r98 <= biasIn_0_r97;
    biasIn_0_r99 <= biasIn_0_r98;
    biasIn_0_r100 <= biasIn_0_r99;
    biasIn_0_r101 <= biasIn_0_r100;
    biasIn_0_r102 <= biasIn_0_r101;
    biasIn_0_r103 <= biasIn_0_r102;
    biasIn_0_r104 <= biasIn_0_r103;
    biasIn_0_r105 <= biasIn_0_r104;
    biasIn_0_r106 <= biasIn_0_r105;
    biasIn_0_r107 <= biasIn_0_r106;
    biasIn_0_r108 <= biasIn_0_r107;
    biasIn_0_r109 <= biasIn_0_r108;
    biasIn_0_r110 <= biasIn_0_r109;
    biasIn_0_r111 <= biasIn_0_r110;
    biasIn_0_r112 <= biasIn_0_r111;
    biasIn_0_r113 <= biasIn_0_r112;
    biasIn_0_r114 <= biasIn_0_r113;
    biasIn_0_r115 <= biasIn_0_r114;
    biasIn_0_r116 <= biasIn_0_r115;
    biasIn_0_r117 <= biasIn_0_r116;
    biasIn_0_r118 <= biasIn_0_r117;
    biasIn_0_r119 <= biasIn_0_r118;
    biasIn_0_r120 <= biasIn_0_r119;
    biasIn_0_r121 <= biasIn_0_r120;
    biasIn_0_r122 <= biasIn_0_r121;
    biasIn_0_r123 <= biasIn_0_r122;
    biasIn_0_r124 <= biasIn_0_r123;
    biasIn_0_r125 <= biasIn_0_r124;
    biasIn_0_r126 <= biasIn_0_r125;
    biasIn_0_r127 <= biasIn_0_r126;
    biasIn_0_r128 <= biasIn_0_r127;
  end
end
////////////////////////////////////////////////////////////////////////////////
// neuron0
////////////////////////////////////////////////////////////////////////////////

neuron neuron0 (
    .biasIn_0(biasIn_0_w0),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w0),
    .reset(reset),
    .tapIn_0(tapIn_0));

////////////////////////////////////////////////////////////////////////////////
// neuron1
////////////////////////////////////////////////////////////////////////////////

neuron neuron1 (
    .biasIn_0(biasIn_0_w1),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w1),
    .reset(reset),
    .tapIn_0(tapIn_1));

////////////////////////////////////////////////////////////////////////////////
// neuron2
////////////////////////////////////////////////////////////////////////////////

neuron neuron2 (
    .biasIn_0(biasIn_0_w2),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w2),
    .reset(reset),
    .tapIn_0(tapIn_2));

////////////////////////////////////////////////////////////////////////////////
// neuron3
////////////////////////////////////////////////////////////////////////////////

neuron neuron3 (
    .biasIn_0(biasIn_0_w3),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w3),
    .reset(reset),
    .tapIn_0(tapIn_3));

////////////////////////////////////////////////////////////////////////////////
// neuron4
////////////////////////////////////////////////////////////////////////////////

neuron neuron4 (
    .biasIn_0(biasIn_0_w4),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w4),
    .reset(reset),
    .tapIn_0(tapIn_4));

////////////////////////////////////////////////////////////////////////////////
// neuron5
////////////////////////////////////////////////////////////////////////////////

neuron neuron5 (
    .biasIn_0(biasIn_0_w5),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w5),
    .reset(reset),
    .tapIn_0(tapIn_5));

////////////////////////////////////////////////////////////////////////////////
// neuron6
////////////////////////////////////////////////////////////////////////////////

neuron neuron6 (
    .biasIn_0(biasIn_0_w6),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w6),
    .reset(reset),
    .tapIn_0(tapIn_6));

////////////////////////////////////////////////////////////////////////////////
// neuron7
////////////////////////////////////////////////////////////////////////////////

neuron neuron7 (
    .biasIn_0(biasIn_0_w7),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w7),
    .reset(reset),
    .tapIn_0(tapIn_7));

////////////////////////////////////////////////////////////////////////////////
// neuron8
////////////////////////////////////////////////////////////////////////////////

neuron neuron8 (
    .biasIn_0(biasIn_0_w8),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w8),
    .reset(reset),
    .tapIn_0(tapIn_8));

////////////////////////////////////////////////////////////////////////////////
// neuron9
////////////////////////////////////////////////////////////////////////////////

neuron neuron9 (
    .biasIn_0(biasIn_0_w9),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w9),
    .reset(reset),
    .tapIn_0(tapIn_9));

////////////////////////////////////////////////////////////////////////////////
// neuron10
////////////////////////////////////////////////////////////////////////////////

neuron neuron10 (
    .biasIn_0(biasIn_0_w10),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w10),
    .reset(reset),
    .tapIn_0(tapIn_10));

////////////////////////////////////////////////////////////////////////////////
// neuron11
////////////////////////////////////////////////////////////////////////////////

neuron neuron11 (
    .biasIn_0(biasIn_0_w11),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w11),
    .reset(reset),
    .tapIn_0(tapIn_11));

////////////////////////////////////////////////////////////////////////////////
// neuron12
////////////////////////////////////////////////////////////////////////////////

neuron neuron12 (
    .biasIn_0(biasIn_0_w12),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w12),
    .reset(reset),
    .tapIn_0(tapIn_12));

////////////////////////////////////////////////////////////////////////////////
// neuron13
////////////////////////////////////////////////////////////////////////////////

neuron neuron13 (
    .biasIn_0(biasIn_0_w13),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w13),
    .reset(reset),
    .tapIn_0(tapIn_13));

////////////////////////////////////////////////////////////////////////////////
// neuron14
////////////////////////////////////////////////////////////////////////////////

neuron neuron14 (
    .biasIn_0(biasIn_0_w14),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w14),
    .reset(reset),
    .tapIn_0(tapIn_14));

////////////////////////////////////////////////////////////////////////////////
// neuron15
////////////////////////////////////////////////////////////////////////////////

neuron neuron15 (
    .biasIn_0(biasIn_0_w15),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w15),
    .reset(reset),
    .tapIn_0(tapIn_15));

////////////////////////////////////////////////////////////////////////////////
// neuron16
////////////////////////////////////////////////////////////////////////////////

neuron neuron16 (
    .biasIn_0(biasIn_0_w16),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w16),
    .reset(reset),
    .tapIn_0(tapIn_16));

////////////////////////////////////////////////////////////////////////////////
// neuron17
////////////////////////////////////////////////////////////////////////////////

neuron neuron17 (
    .biasIn_0(biasIn_0_w17),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w17),
    .reset(reset),
    .tapIn_0(tapIn_17));

////////////////////////////////////////////////////////////////////////////////
// neuron18
////////////////////////////////////////////////////////////////////////////////

neuron neuron18 (
    .biasIn_0(biasIn_0_w18),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w18),
    .reset(reset),
    .tapIn_0(tapIn_18));

////////////////////////////////////////////////////////////////////////////////
// neuron19
////////////////////////////////////////////////////////////////////////////////

neuron neuron19 (
    .biasIn_0(biasIn_0_w19),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w19),
    .reset(reset),
    .tapIn_0(tapIn_19));

////////////////////////////////////////////////////////////////////////////////
// neuron20
////////////////////////////////////////////////////////////////////////////////

neuron neuron20 (
    .biasIn_0(biasIn_0_w20),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w20),
    .reset(reset),
    .tapIn_0(tapIn_20));

////////////////////////////////////////////////////////////////////////////////
// neuron21
////////////////////////////////////////////////////////////////////////////////

neuron neuron21 (
    .biasIn_0(biasIn_0_w21),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w21),
    .reset(reset),
    .tapIn_0(tapIn_21));

////////////////////////////////////////////////////////////////////////////////
// neuron22
////////////////////////////////////////////////////////////////////////////////

neuron neuron22 (
    .biasIn_0(biasIn_0_w22),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w22),
    .reset(reset),
    .tapIn_0(tapIn_22));

////////////////////////////////////////////////////////////////////////////////
// neuron23
////////////////////////////////////////////////////////////////////////////////

neuron neuron23 (
    .biasIn_0(biasIn_0_w23),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w23),
    .reset(reset),
    .tapIn_0(tapIn_23));

////////////////////////////////////////////////////////////////////////////////
// neuron24
////////////////////////////////////////////////////////////////////////////////

neuron neuron24 (
    .biasIn_0(biasIn_0_w24),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w24),
    .reset(reset),
    .tapIn_0(tapIn_24));

////////////////////////////////////////////////////////////////////////////////
// neuron25
////////////////////////////////////////////////////////////////////////////////

neuron neuron25 (
    .biasIn_0(biasIn_0_w25),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w25),
    .reset(reset),
    .tapIn_0(tapIn_25));

////////////////////////////////////////////////////////////////////////////////
// neuron26
////////////////////////////////////////////////////////////////////////////////

neuron neuron26 (
    .biasIn_0(biasIn_0_w26),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w26),
    .reset(reset),
    .tapIn_0(tapIn_26));

////////////////////////////////////////////////////////////////////////////////
// neuron27
////////////////////////////////////////////////////////////////////////////////

neuron neuron27 (
    .biasIn_0(biasIn_0_w27),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w27),
    .reset(reset),
    .tapIn_0(tapIn_27));

////////////////////////////////////////////////////////////////////////////////
// neuron28
////////////////////////////////////////////////////////////////////////////////

neuron neuron28 (
    .biasIn_0(biasIn_0_w28),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w28),
    .reset(reset),
    .tapIn_0(tapIn_28));

////////////////////////////////////////////////////////////////////////////////
// neuron29
////////////////////////////////////////////////////////////////////////////////

neuron neuron29 (
    .biasIn_0(biasIn_0_w29),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w29),
    .reset(reset),
    .tapIn_0(tapIn_29));

////////////////////////////////////////////////////////////////////////////////
// neuron30
////////////////////////////////////////////////////////////////////////////////

neuron neuron30 (
    .biasIn_0(biasIn_0_w30),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w30),
    .reset(reset),
    .tapIn_0(tapIn_30));

////////////////////////////////////////////////////////////////////////////////
// neuron31
////////////////////////////////////////////////////////////////////////////////

neuron neuron31 (
    .biasIn_0(biasIn_0_w31),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w31),
    .reset(reset),
    .tapIn_0(tapIn_31));

////////////////////////////////////////////////////////////////////////////////
// neuron32
////////////////////////////////////////////////////////////////////////////////

neuron neuron32 (
    .biasIn_0(biasIn_0_w32),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w32),
    .reset(reset),
    .tapIn_0(tapIn_32));

////////////////////////////////////////////////////////////////////////////////
// neuron33
////////////////////////////////////////////////////////////////////////////////

neuron neuron33 (
    .biasIn_0(biasIn_0_w33),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w33),
    .reset(reset),
    .tapIn_0(tapIn_33));

////////////////////////////////////////////////////////////////////////////////
// neuron34
////////////////////////////////////////////////////////////////////////////////

neuron neuron34 (
    .biasIn_0(biasIn_0_w34),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w34),
    .reset(reset),
    .tapIn_0(tapIn_34));

////////////////////////////////////////////////////////////////////////////////
// neuron35
////////////////////////////////////////////////////////////////////////////////

neuron neuron35 (
    .biasIn_0(biasIn_0_w35),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w35),
    .reset(reset),
    .tapIn_0(tapIn_35));

////////////////////////////////////////////////////////////////////////////////
// neuron36
////////////////////////////////////////////////////////////////////////////////

neuron neuron36 (
    .biasIn_0(biasIn_0_w36),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w36),
    .reset(reset),
    .tapIn_0(tapIn_36));

////////////////////////////////////////////////////////////////////////////////
// neuron37
////////////////////////////////////////////////////////////////////////////////

neuron neuron37 (
    .biasIn_0(biasIn_0_w37),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w37),
    .reset(reset),
    .tapIn_0(tapIn_37));

////////////////////////////////////////////////////////////////////////////////
// neuron38
////////////////////////////////////////////////////////////////////////////////

neuron neuron38 (
    .biasIn_0(biasIn_0_w38),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w38),
    .reset(reset),
    .tapIn_0(tapIn_38));

////////////////////////////////////////////////////////////////////////////////
// neuron39
////////////////////////////////////////////////////////////////////////////////

neuron neuron39 (
    .biasIn_0(biasIn_0_w39),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w39),
    .reset(reset),
    .tapIn_0(tapIn_39));

////////////////////////////////////////////////////////////////////////////////
// neuron40
////////////////////////////////////////////////////////////////////////////////

neuron neuron40 (
    .biasIn_0(biasIn_0_w40),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w40),
    .reset(reset),
    .tapIn_0(tapIn_40));

////////////////////////////////////////////////////////////////////////////////
// neuron41
////////////////////////////////////////////////////////////////////////////////

neuron neuron41 (
    .biasIn_0(biasIn_0_w41),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w41),
    .reset(reset),
    .tapIn_0(tapIn_41));

////////////////////////////////////////////////////////////////////////////////
// neuron42
////////////////////////////////////////////////////////////////////////////////

neuron neuron42 (
    .biasIn_0(biasIn_0_w42),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w42),
    .reset(reset),
    .tapIn_0(tapIn_42));

////////////////////////////////////////////////////////////////////////////////
// neuron43
////////////////////////////////////////////////////////////////////////////////

neuron neuron43 (
    .biasIn_0(biasIn_0_w43),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w43),
    .reset(reset),
    .tapIn_0(tapIn_43));

////////////////////////////////////////////////////////////////////////////////
// neuron44
////////////////////////////////////////////////////////////////////////////////

neuron neuron44 (
    .biasIn_0(biasIn_0_w44),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w44),
    .reset(reset),
    .tapIn_0(tapIn_44));

////////////////////////////////////////////////////////////////////////////////
// neuron45
////////////////////////////////////////////////////////////////////////////////

neuron neuron45 (
    .biasIn_0(biasIn_0_w45),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w45),
    .reset(reset),
    .tapIn_0(tapIn_45));

////////////////////////////////////////////////////////////////////////////////
// neuron46
////////////////////////////////////////////////////////////////////////////////

neuron neuron46 (
    .biasIn_0(biasIn_0_w46),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w46),
    .reset(reset),
    .tapIn_0(tapIn_46));

////////////////////////////////////////////////////////////////////////////////
// neuron47
////////////////////////////////////////////////////////////////////////////////

neuron neuron47 (
    .biasIn_0(biasIn_0_w47),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w47),
    .reset(reset),
    .tapIn_0(tapIn_47));

////////////////////////////////////////////////////////////////////////////////
// neuron48
////////////////////////////////////////////////////////////////////////////////

neuron neuron48 (
    .biasIn_0(biasIn_0_w48),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w48),
    .reset(reset),
    .tapIn_0(tapIn_48));

////////////////////////////////////////////////////////////////////////////////
// neuron49
////////////////////////////////////////////////////////////////////////////////

neuron neuron49 (
    .biasIn_0(biasIn_0_w49),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w49),
    .reset(reset),
    .tapIn_0(tapIn_49));

////////////////////////////////////////////////////////////////////////////////
// neuron50
////////////////////////////////////////////////////////////////////////////////

neuron neuron50 (
    .biasIn_0(biasIn_0_w50),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w50),
    .reset(reset),
    .tapIn_0(tapIn_50));

////////////////////////////////////////////////////////////////////////////////
// neuron51
////////////////////////////////////////////////////////////////////////////////

neuron neuron51 (
    .biasIn_0(biasIn_0_w51),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w51),
    .reset(reset),
    .tapIn_0(tapIn_51));

////////////////////////////////////////////////////////////////////////////////
// neuron52
////////////////////////////////////////////////////////////////////////////////

neuron neuron52 (
    .biasIn_0(biasIn_0_w52),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w52),
    .reset(reset),
    .tapIn_0(tapIn_52));

////////////////////////////////////////////////////////////////////////////////
// neuron53
////////////////////////////////////////////////////////////////////////////////

neuron neuron53 (
    .biasIn_0(biasIn_0_w53),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w53),
    .reset(reset),
    .tapIn_0(tapIn_53));

////////////////////////////////////////////////////////////////////////////////
// neuron54
////////////////////////////////////////////////////////////////////////////////

neuron neuron54 (
    .biasIn_0(biasIn_0_w54),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w54),
    .reset(reset),
    .tapIn_0(tapIn_54));

////////////////////////////////////////////////////////////////////////////////
// neuron55
////////////////////////////////////////////////////////////////////////////////

neuron neuron55 (
    .biasIn_0(biasIn_0_w55),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w55),
    .reset(reset),
    .tapIn_0(tapIn_55));

////////////////////////////////////////////////////////////////////////////////
// neuron56
////////////////////////////////////////////////////////////////////////////////

neuron neuron56 (
    .biasIn_0(biasIn_0_w56),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w56),
    .reset(reset),
    .tapIn_0(tapIn_56));

////////////////////////////////////////////////////////////////////////////////
// neuron57
////////////////////////////////////////////////////////////////////////////////

neuron neuron57 (
    .biasIn_0(biasIn_0_w57),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w57),
    .reset(reset),
    .tapIn_0(tapIn_57));

////////////////////////////////////////////////////////////////////////////////
// neuron58
////////////////////////////////////////////////////////////////////////////////

neuron neuron58 (
    .biasIn_0(biasIn_0_w58),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w58),
    .reset(reset),
    .tapIn_0(tapIn_58));

////////////////////////////////////////////////////////////////////////////////
// neuron59
////////////////////////////////////////////////////////////////////////////////

neuron neuron59 (
    .biasIn_0(biasIn_0_w59),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w59),
    .reset(reset),
    .tapIn_0(tapIn_59));

////////////////////////////////////////////////////////////////////////////////
// neuron60
////////////////////////////////////////////////////////////////////////////////

neuron neuron60 (
    .biasIn_0(biasIn_0_w60),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w60),
    .reset(reset),
    .tapIn_0(tapIn_60));

////////////////////////////////////////////////////////////////////////////////
// neuron61
////////////////////////////////////////////////////////////////////////////////

neuron neuron61 (
    .biasIn_0(biasIn_0_w61),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w61),
    .reset(reset),
    .tapIn_0(tapIn_61));

////////////////////////////////////////////////////////////////////////////////
// neuron62
////////////////////////////////////////////////////////////////////////////////

neuron neuron62 (
    .biasIn_0(biasIn_0_w62),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w62),
    .reset(reset),
    .tapIn_0(tapIn_62));

////////////////////////////////////////////////////////////////////////////////
// neuron63
////////////////////////////////////////////////////////////////////////////////

neuron neuron63 (
    .biasIn_0(biasIn_0_w63),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w63),
    .reset(reset),
    .tapIn_0(tapIn_63));

////////////////////////////////////////////////////////////////////////////////
// neuron64
////////////////////////////////////////////////////////////////////////////////

neuron neuron64 (
    .biasIn_0(biasIn_0_w64),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w64),
    .reset(reset),
    .tapIn_0(tapIn_64));

////////////////////////////////////////////////////////////////////////////////
// neuron65
////////////////////////////////////////////////////////////////////////////////

neuron neuron65 (
    .biasIn_0(biasIn_0_w65),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w65),
    .reset(reset),
    .tapIn_0(tapIn_65));

////////////////////////////////////////////////////////////////////////////////
// neuron66
////////////////////////////////////////////////////////////////////////////////

neuron neuron66 (
    .biasIn_0(biasIn_0_w66),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w66),
    .reset(reset),
    .tapIn_0(tapIn_66));

////////////////////////////////////////////////////////////////////////////////
// neuron67
////////////////////////////////////////////////////////////////////////////////

neuron neuron67 (
    .biasIn_0(biasIn_0_w67),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w67),
    .reset(reset),
    .tapIn_0(tapIn_67));

////////////////////////////////////////////////////////////////////////////////
// neuron68
////////////////////////////////////////////////////////////////////////////////

neuron neuron68 (
    .biasIn_0(biasIn_0_w68),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w68),
    .reset(reset),
    .tapIn_0(tapIn_68));

////////////////////////////////////////////////////////////////////////////////
// neuron69
////////////////////////////////////////////////////////////////////////////////

neuron neuron69 (
    .biasIn_0(biasIn_0_w69),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w69),
    .reset(reset),
    .tapIn_0(tapIn_69));

////////////////////////////////////////////////////////////////////////////////
// neuron70
////////////////////////////////////////////////////////////////////////////////

neuron neuron70 (
    .biasIn_0(biasIn_0_w70),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w70),
    .reset(reset),
    .tapIn_0(tapIn_70));

////////////////////////////////////////////////////////////////////////////////
// neuron71
////////////////////////////////////////////////////////////////////////////////

neuron neuron71 (
    .biasIn_0(biasIn_0_w71),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w71),
    .reset(reset),
    .tapIn_0(tapIn_71));

////////////////////////////////////////////////////////////////////////////////
// neuron72
////////////////////////////////////////////////////////////////////////////////

neuron neuron72 (
    .biasIn_0(biasIn_0_w72),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w72),
    .reset(reset),
    .tapIn_0(tapIn_72));

////////////////////////////////////////////////////////////////////////////////
// neuron73
////////////////////////////////////////////////////////////////////////////////

neuron neuron73 (
    .biasIn_0(biasIn_0_w73),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w73),
    .reset(reset),
    .tapIn_0(tapIn_73));

////////////////////////////////////////////////////////////////////////////////
// neuron74
////////////////////////////////////////////////////////////////////////////////

neuron neuron74 (
    .biasIn_0(biasIn_0_w74),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w74),
    .reset(reset),
    .tapIn_0(tapIn_74));

////////////////////////////////////////////////////////////////////////////////
// neuron75
////////////////////////////////////////////////////////////////////////////////

neuron neuron75 (
    .biasIn_0(biasIn_0_w75),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w75),
    .reset(reset),
    .tapIn_0(tapIn_75));

////////////////////////////////////////////////////////////////////////////////
// neuron76
////////////////////////////////////////////////////////////////////////////////

neuron neuron76 (
    .biasIn_0(biasIn_0_w76),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w76),
    .reset(reset),
    .tapIn_0(tapIn_76));

////////////////////////////////////////////////////////////////////////////////
// neuron77
////////////////////////////////////////////////////////////////////////////////

neuron neuron77 (
    .biasIn_0(biasIn_0_w77),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w77),
    .reset(reset),
    .tapIn_0(tapIn_77));

////////////////////////////////////////////////////////////////////////////////
// neuron78
////////////////////////////////////////////////////////////////////////////////

neuron neuron78 (
    .biasIn_0(biasIn_0_w78),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w78),
    .reset(reset),
    .tapIn_0(tapIn_78));

////////////////////////////////////////////////////////////////////////////////
// neuron79
////////////////////////////////////////////////////////////////////////////////

neuron neuron79 (
    .biasIn_0(biasIn_0_w79),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w79),
    .reset(reset),
    .tapIn_0(tapIn_79));

////////////////////////////////////////////////////////////////////////////////
// neuron80
////////////////////////////////////////////////////////////////////////////////

neuron neuron80 (
    .biasIn_0(biasIn_0_w80),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w80),
    .reset(reset),
    .tapIn_0(tapIn_80));

////////////////////////////////////////////////////////////////////////////////
// neuron81
////////////////////////////////////////////////////////////////////////////////

neuron neuron81 (
    .biasIn_0(biasIn_0_w81),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w81),
    .reset(reset),
    .tapIn_0(tapIn_81));

////////////////////////////////////////////////////////////////////////////////
// neuron82
////////////////////////////////////////////////////////////////////////////////

neuron neuron82 (
    .biasIn_0(biasIn_0_w82),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w82),
    .reset(reset),
    .tapIn_0(tapIn_82));

////////////////////////////////////////////////////////////////////////////////
// neuron83
////////////////////////////////////////////////////////////////////////////////

neuron neuron83 (
    .biasIn_0(biasIn_0_w83),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w83),
    .reset(reset),
    .tapIn_0(tapIn_83));

////////////////////////////////////////////////////////////////////////////////
// neuron84
////////////////////////////////////////////////////////////////////////////////

neuron neuron84 (
    .biasIn_0(biasIn_0_w84),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w84),
    .reset(reset),
    .tapIn_0(tapIn_84));

////////////////////////////////////////////////////////////////////////////////
// neuron85
////////////////////////////////////////////////////////////////////////////////

neuron neuron85 (
    .biasIn_0(biasIn_0_w85),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w85),
    .reset(reset),
    .tapIn_0(tapIn_85));

////////////////////////////////////////////////////////////////////////////////
// neuron86
////////////////////////////////////////////////////////////////////////////////

neuron neuron86 (
    .biasIn_0(biasIn_0_w86),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w86),
    .reset(reset),
    .tapIn_0(tapIn_86));

////////////////////////////////////////////////////////////////////////////////
// neuron87
////////////////////////////////////////////////////////////////////////////////

neuron neuron87 (
    .biasIn_0(biasIn_0_w87),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w87),
    .reset(reset),
    .tapIn_0(tapIn_87));

////////////////////////////////////////////////////////////////////////////////
// neuron88
////////////////////////////////////////////////////////////////////////////////

neuron neuron88 (
    .biasIn_0(biasIn_0_w88),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w88),
    .reset(reset),
    .tapIn_0(tapIn_88));

////////////////////////////////////////////////////////////////////////////////
// neuron89
////////////////////////////////////////////////////////////////////////////////

neuron neuron89 (
    .biasIn_0(biasIn_0_w89),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w89),
    .reset(reset),
    .tapIn_0(tapIn_89));

////////////////////////////////////////////////////////////////////////////////
// neuron90
////////////////////////////////////////////////////////////////////////////////

neuron neuron90 (
    .biasIn_0(biasIn_0_w90),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w90),
    .reset(reset),
    .tapIn_0(tapIn_90));

////////////////////////////////////////////////////////////////////////////////
// neuron91
////////////////////////////////////////////////////////////////////////////////

neuron neuron91 (
    .biasIn_0(biasIn_0_w91),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w91),
    .reset(reset),
    .tapIn_0(tapIn_91));

////////////////////////////////////////////////////////////////////////////////
// neuron92
////////////////////////////////////////////////////////////////////////////////

neuron neuron92 (
    .biasIn_0(biasIn_0_w92),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w92),
    .reset(reset),
    .tapIn_0(tapIn_92));

////////////////////////////////////////////////////////////////////////////////
// neuron93
////////////////////////////////////////////////////////////////////////////////

neuron neuron93 (
    .biasIn_0(biasIn_0_w93),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w93),
    .reset(reset),
    .tapIn_0(tapIn_93));

////////////////////////////////////////////////////////////////////////////////
// neuron94
////////////////////////////////////////////////////////////////////////////////

neuron neuron94 (
    .biasIn_0(biasIn_0_w94),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w94),
    .reset(reset),
    .tapIn_0(tapIn_94));

////////////////////////////////////////////////////////////////////////////////
// neuron95
////////////////////////////////////////////////////////////////////////////////

neuron neuron95 (
    .biasIn_0(biasIn_0_w95),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w95),
    .reset(reset),
    .tapIn_0(tapIn_95));

////////////////////////////////////////////////////////////////////////////////
// neuron96
////////////////////////////////////////////////////////////////////////////////

neuron neuron96 (
    .biasIn_0(biasIn_0_w96),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w96),
    .reset(reset),
    .tapIn_0(tapIn_96));

////////////////////////////////////////////////////////////////////////////////
// neuron97
////////////////////////////////////////////////////////////////////////////////

neuron neuron97 (
    .biasIn_0(biasIn_0_w97),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w97),
    .reset(reset),
    .tapIn_0(tapIn_97));

////////////////////////////////////////////////////////////////////////////////
// neuron98
////////////////////////////////////////////////////////////////////////////////

neuron neuron98 (
    .biasIn_0(biasIn_0_w98),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w98),
    .reset(reset),
    .tapIn_0(tapIn_98));

////////////////////////////////////////////////////////////////////////////////
// neuron99
////////////////////////////////////////////////////////////////////////////////

neuron neuron99 (
    .biasIn_0(biasIn_0_w99),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w99),
    .reset(reset),
    .tapIn_0(tapIn_99));

////////////////////////////////////////////////////////////////////////////////
// neuron100
////////////////////////////////////////////////////////////////////////////////

neuron neuron100 (
    .biasIn_0(biasIn_0_w100),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w100),
    .reset(reset),
    .tapIn_0(tapIn_100));

////////////////////////////////////////////////////////////////////////////////
// neuron101
////////////////////////////////////////////////////////////////////////////////

neuron neuron101 (
    .biasIn_0(biasIn_0_w101),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w101),
    .reset(reset),
    .tapIn_0(tapIn_101));

////////////////////////////////////////////////////////////////////////////////
// neuron102
////////////////////////////////////////////////////////////////////////////////

neuron neuron102 (
    .biasIn_0(biasIn_0_w102),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w102),
    .reset(reset),
    .tapIn_0(tapIn_102));

////////////////////////////////////////////////////////////////////////////////
// neuron103
////////////////////////////////////////////////////////////////////////////////

neuron neuron103 (
    .biasIn_0(biasIn_0_w103),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w103),
    .reset(reset),
    .tapIn_0(tapIn_103));

////////////////////////////////////////////////////////////////////////////////
// neuron104
////////////////////////////////////////////////////////////////////////////////

neuron neuron104 (
    .biasIn_0(biasIn_0_w104),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w104),
    .reset(reset),
    .tapIn_0(tapIn_104));

////////////////////////////////////////////////////////////////////////////////
// neuron105
////////////////////////////////////////////////////////////////////////////////

neuron neuron105 (
    .biasIn_0(biasIn_0_w105),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w105),
    .reset(reset),
    .tapIn_0(tapIn_105));

////////////////////////////////////////////////////////////////////////////////
// neuron106
////////////////////////////////////////////////////////////////////////////////

neuron neuron106 (
    .biasIn_0(biasIn_0_w106),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w106),
    .reset(reset),
    .tapIn_0(tapIn_106));

////////////////////////////////////////////////////////////////////////////////
// neuron107
////////////////////////////////////////////////////////////////////////////////

neuron neuron107 (
    .biasIn_0(biasIn_0_w107),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w107),
    .reset(reset),
    .tapIn_0(tapIn_107));

////////////////////////////////////////////////////////////////////////////////
// neuron108
////////////////////////////////////////////////////////////////////////////////

neuron neuron108 (
    .biasIn_0(biasIn_0_w108),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w108),
    .reset(reset),
    .tapIn_0(tapIn_108));

////////////////////////////////////////////////////////////////////////////////
// neuron109
////////////////////////////////////////////////////////////////////////////////

neuron neuron109 (
    .biasIn_0(biasIn_0_w109),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w109),
    .reset(reset),
    .tapIn_0(tapIn_109));

////////////////////////////////////////////////////////////////////////////////
// neuron110
////////////////////////////////////////////////////////////////////////////////

neuron neuron110 (
    .biasIn_0(biasIn_0_w110),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w110),
    .reset(reset),
    .tapIn_0(tapIn_110));

////////////////////////////////////////////////////////////////////////////////
// neuron111
////////////////////////////////////////////////////////////////////////////////

neuron neuron111 (
    .biasIn_0(biasIn_0_w111),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w111),
    .reset(reset),
    .tapIn_0(tapIn_111));

////////////////////////////////////////////////////////////////////////////////
// neuron112
////////////////////////////////////////////////////////////////////////////////

neuron neuron112 (
    .biasIn_0(biasIn_0_w112),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w112),
    .reset(reset),
    .tapIn_0(tapIn_112));

////////////////////////////////////////////////////////////////////////////////
// neuron113
////////////////////////////////////////////////////////////////////////////////

neuron neuron113 (
    .biasIn_0(biasIn_0_w113),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w113),
    .reset(reset),
    .tapIn_0(tapIn_113));

////////////////////////////////////////////////////////////////////////////////
// neuron114
////////////////////////////////////////////////////////////////////////////////

neuron neuron114 (
    .biasIn_0(biasIn_0_w114),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w114),
    .reset(reset),
    .tapIn_0(tapIn_114));

////////////////////////////////////////////////////////////////////////////////
// neuron115
////////////////////////////////////////////////////////////////////////////////

neuron neuron115 (
    .biasIn_0(biasIn_0_w115),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w115),
    .reset(reset),
    .tapIn_0(tapIn_115));

////////////////////////////////////////////////////////////////////////////////
// neuron116
////////////////////////////////////////////////////////////////////////////////

neuron neuron116 (
    .biasIn_0(biasIn_0_w116),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w116),
    .reset(reset),
    .tapIn_0(tapIn_116));

////////////////////////////////////////////////////////////////////////////////
// neuron117
////////////////////////////////////////////////////////////////////////////////

neuron neuron117 (
    .biasIn_0(biasIn_0_w117),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w117),
    .reset(reset),
    .tapIn_0(tapIn_117));

////////////////////////////////////////////////////////////////////////////////
// neuron118
////////////////////////////////////////////////////////////////////////////////

neuron neuron118 (
    .biasIn_0(biasIn_0_w118),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w118),
    .reset(reset),
    .tapIn_0(tapIn_118));

////////////////////////////////////////////////////////////////////////////////
// neuron119
////////////////////////////////////////////////////////////////////////////////

neuron neuron119 (
    .biasIn_0(biasIn_0_w119),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w119),
    .reset(reset),
    .tapIn_0(tapIn_119));

////////////////////////////////////////////////////////////////////////////////
// neuron120
////////////////////////////////////////////////////////////////////////////////

neuron neuron120 (
    .biasIn_0(biasIn_0_w120),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w120),
    .reset(reset),
    .tapIn_0(tapIn_120));

////////////////////////////////////////////////////////////////////////////////
// neuron121
////////////////////////////////////////////////////////////////////////////////

neuron neuron121 (
    .biasIn_0(biasIn_0_w121),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w121),
    .reset(reset),
    .tapIn_0(tapIn_121));

////////////////////////////////////////////////////////////////////////////////
// neuron122
////////////////////////////////////////////////////////////////////////////////

neuron neuron122 (
    .biasIn_0(biasIn_0_w122),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w122),
    .reset(reset),
    .tapIn_0(tapIn_122));

////////////////////////////////////////////////////////////////////////////////
// neuron123
////////////////////////////////////////////////////////////////////////////////

neuron neuron123 (
    .biasIn_0(biasIn_0_w123),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w123),
    .reset(reset),
    .tapIn_0(tapIn_123));

////////////////////////////////////////////////////////////////////////////////
// neuron124
////////////////////////////////////////////////////////////////////////////////

neuron neuron124 (
    .biasIn_0(biasIn_0_w124),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w124),
    .reset(reset),
    .tapIn_0(tapIn_124));

////////////////////////////////////////////////////////////////////////////////
// neuron125
////////////////////////////////////////////////////////////////////////////////

neuron neuron125 (
    .biasIn_0(biasIn_0_w125),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w125),
    .reset(reset),
    .tapIn_0(tapIn_125));

////////////////////////////////////////////////////////////////////////////////
// neuron126
////////////////////////////////////////////////////////////////////////////////

neuron neuron126 (
    .biasIn_0(biasIn_0_w126),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w126),
    .reset(reset),
    .tapIn_0(tapIn_126));

////////////////////////////////////////////////////////////////////////////////
// neuron127
////////////////////////////////////////////////////////////////////////////////

neuron neuron127 (
    .biasIn_0(biasIn_0_w127),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOut_0(wireOut_w127),
    .reset(reset),
    .tapIn_0(tapIn_127));

////////////////////////////////////////////////////////////////////////////////
// sigmoid
////////////////////////////////////////////////////////////////////////////////

sigmoid sigmoid (
    .clk(clk),
    .dataOutPre_0(outLine_w0),
    .dataOut_0(dataOut_0),
    .reset(reset));


// Delay the Input Valid
always @(posedge clk) begin
  if (reset) begin
    valid0 <= 'd0;
    valid1 <= 'd0;
  end
  else begin
    valid0 <= valid;
    valid1 <= valid0;
  end
end

// Select the inputs to the Neuron

assign biasIn_0_w0 = valid0 ? biasIn_0_r127 : wireOut_w0;
assign biasIn_0_w1 = valid0 ? biasIn_0_r126 : wireOut_w1;
assign biasIn_0_w2 = valid0 ? biasIn_0_r125 : wireOut_w2;
assign biasIn_0_w3 = valid0 ? biasIn_0_r124 : wireOut_w3;
assign biasIn_0_w4 = valid0 ? biasIn_0_r123 : wireOut_w4;
assign biasIn_0_w5 = valid0 ? biasIn_0_r122 : wireOut_w5;
assign biasIn_0_w6 = valid0 ? biasIn_0_r121 : wireOut_w6;
assign biasIn_0_w7 = valid0 ? biasIn_0_r120 : wireOut_w7;
assign biasIn_0_w8 = valid0 ? biasIn_0_r119 : wireOut_w8;
assign biasIn_0_w9 = valid0 ? biasIn_0_r118 : wireOut_w9;
assign biasIn_0_w10 = valid0 ? biasIn_0_r117 : wireOut_w10;
assign biasIn_0_w11 = valid0 ? biasIn_0_r116 : wireOut_w11;
assign biasIn_0_w12 = valid0 ? biasIn_0_r115 : wireOut_w12;
assign biasIn_0_w13 = valid0 ? biasIn_0_r114 : wireOut_w13;
assign biasIn_0_w14 = valid0 ? biasIn_0_r113 : wireOut_w14;
assign biasIn_0_w15 = valid0 ? biasIn_0_r112 : wireOut_w15;
assign biasIn_0_w16 = valid0 ? biasIn_0_r111 : wireOut_w16;
assign biasIn_0_w17 = valid0 ? biasIn_0_r110 : wireOut_w17;
assign biasIn_0_w18 = valid0 ? biasIn_0_r109 : wireOut_w18;
assign biasIn_0_w19 = valid0 ? biasIn_0_r108 : wireOut_w19;
assign biasIn_0_w20 = valid0 ? biasIn_0_r107 : wireOut_w20;
assign biasIn_0_w21 = valid0 ? biasIn_0_r106 : wireOut_w21;
assign biasIn_0_w22 = valid0 ? biasIn_0_r105 : wireOut_w22;
assign biasIn_0_w23 = valid0 ? biasIn_0_r104 : wireOut_w23;
assign biasIn_0_w24 = valid0 ? biasIn_0_r103 : wireOut_w24;
assign biasIn_0_w25 = valid0 ? biasIn_0_r102 : wireOut_w25;
assign biasIn_0_w26 = valid0 ? biasIn_0_r101 : wireOut_w26;
assign biasIn_0_w27 = valid0 ? biasIn_0_r100 : wireOut_w27;
assign biasIn_0_w28 = valid0 ? biasIn_0_r99 : wireOut_w28;
assign biasIn_0_w29 = valid0 ? biasIn_0_r98 : wireOut_w29;
assign biasIn_0_w30 = valid0 ? biasIn_0_r97 : wireOut_w30;
assign biasIn_0_w31 = valid0 ? biasIn_0_r96 : wireOut_w31;
assign biasIn_0_w32 = valid0 ? biasIn_0_r95 : wireOut_w32;
assign biasIn_0_w33 = valid0 ? biasIn_0_r94 : wireOut_w33;
assign biasIn_0_w34 = valid0 ? biasIn_0_r93 : wireOut_w34;
assign biasIn_0_w35 = valid0 ? biasIn_0_r92 : wireOut_w35;
assign biasIn_0_w36 = valid0 ? biasIn_0_r91 : wireOut_w36;
assign biasIn_0_w37 = valid0 ? biasIn_0_r90 : wireOut_w37;
assign biasIn_0_w38 = valid0 ? biasIn_0_r89 : wireOut_w38;
assign biasIn_0_w39 = valid0 ? biasIn_0_r88 : wireOut_w39;
assign biasIn_0_w40 = valid0 ? biasIn_0_r87 : wireOut_w40;
assign biasIn_0_w41 = valid0 ? biasIn_0_r86 : wireOut_w41;
assign biasIn_0_w42 = valid0 ? biasIn_0_r85 : wireOut_w42;
assign biasIn_0_w43 = valid0 ? biasIn_0_r84 : wireOut_w43;
assign biasIn_0_w44 = valid0 ? biasIn_0_r83 : wireOut_w44;
assign biasIn_0_w45 = valid0 ? biasIn_0_r82 : wireOut_w45;
assign biasIn_0_w46 = valid0 ? biasIn_0_r81 : wireOut_w46;
assign biasIn_0_w47 = valid0 ? biasIn_0_r80 : wireOut_w47;
assign biasIn_0_w48 = valid0 ? biasIn_0_r79 : wireOut_w48;
assign biasIn_0_w49 = valid0 ? biasIn_0_r78 : wireOut_w49;
assign biasIn_0_w50 = valid0 ? biasIn_0_r77 : wireOut_w50;
assign biasIn_0_w51 = valid0 ? biasIn_0_r76 : wireOut_w51;
assign biasIn_0_w52 = valid0 ? biasIn_0_r75 : wireOut_w52;
assign biasIn_0_w53 = valid0 ? biasIn_0_r74 : wireOut_w53;
assign biasIn_0_w54 = valid0 ? biasIn_0_r73 : wireOut_w54;
assign biasIn_0_w55 = valid0 ? biasIn_0_r72 : wireOut_w55;
assign biasIn_0_w56 = valid0 ? biasIn_0_r71 : wireOut_w56;
assign biasIn_0_w57 = valid0 ? biasIn_0_r70 : wireOut_w57;
assign biasIn_0_w58 = valid0 ? biasIn_0_r69 : wireOut_w58;
assign biasIn_0_w59 = valid0 ? biasIn_0_r68 : wireOut_w59;
assign biasIn_0_w60 = valid0 ? biasIn_0_r67 : wireOut_w60;
assign biasIn_0_w61 = valid0 ? biasIn_0_r66 : wireOut_w61;
assign biasIn_0_w62 = valid0 ? biasIn_0_r65 : wireOut_w62;
assign biasIn_0_w63 = valid0 ? biasIn_0_r64 : wireOut_w63;
assign biasIn_0_w64 = valid0 ? biasIn_0_r63 : wireOut_w64;
assign biasIn_0_w65 = valid0 ? biasIn_0_r62 : wireOut_w65;
assign biasIn_0_w66 = valid0 ? biasIn_0_r61 : wireOut_w66;
assign biasIn_0_w67 = valid0 ? biasIn_0_r60 : wireOut_w67;
assign biasIn_0_w68 = valid0 ? biasIn_0_r59 : wireOut_w68;
assign biasIn_0_w69 = valid0 ? biasIn_0_r58 : wireOut_w69;
assign biasIn_0_w70 = valid0 ? biasIn_0_r57 : wireOut_w70;
assign biasIn_0_w71 = valid0 ? biasIn_0_r56 : wireOut_w71;
assign biasIn_0_w72 = valid0 ? biasIn_0_r55 : wireOut_w72;
assign biasIn_0_w73 = valid0 ? biasIn_0_r54 : wireOut_w73;
assign biasIn_0_w74 = valid0 ? biasIn_0_r53 : wireOut_w74;
assign biasIn_0_w75 = valid0 ? biasIn_0_r52 : wireOut_w75;
assign biasIn_0_w76 = valid0 ? biasIn_0_r51 : wireOut_w76;
assign biasIn_0_w77 = valid0 ? biasIn_0_r50 : wireOut_w77;
assign biasIn_0_w78 = valid0 ? biasIn_0_r49 : wireOut_w78;
assign biasIn_0_w79 = valid0 ? biasIn_0_r48 : wireOut_w79;
assign biasIn_0_w80 = valid0 ? biasIn_0_r47 : wireOut_w80;
assign biasIn_0_w81 = valid0 ? biasIn_0_r46 : wireOut_w81;
assign biasIn_0_w82 = valid0 ? biasIn_0_r45 : wireOut_w82;
assign biasIn_0_w83 = valid0 ? biasIn_0_r44 : wireOut_w83;
assign biasIn_0_w84 = valid0 ? biasIn_0_r43 : wireOut_w84;
assign biasIn_0_w85 = valid0 ? biasIn_0_r42 : wireOut_w85;
assign biasIn_0_w86 = valid0 ? biasIn_0_r41 : wireOut_w86;
assign biasIn_0_w87 = valid0 ? biasIn_0_r40 : wireOut_w87;
assign biasIn_0_w88 = valid0 ? biasIn_0_r39 : wireOut_w88;
assign biasIn_0_w89 = valid0 ? biasIn_0_r38 : wireOut_w89;
assign biasIn_0_w90 = valid0 ? biasIn_0_r37 : wireOut_w90;
assign biasIn_0_w91 = valid0 ? biasIn_0_r36 : wireOut_w91;
assign biasIn_0_w92 = valid0 ? biasIn_0_r35 : wireOut_w92;
assign biasIn_0_w93 = valid0 ? biasIn_0_r34 : wireOut_w93;
assign biasIn_0_w94 = valid0 ? biasIn_0_r33 : wireOut_w94;
assign biasIn_0_w95 = valid0 ? biasIn_0_r32 : wireOut_w95;
assign biasIn_0_w96 = valid0 ? biasIn_0_r31 : wireOut_w96;
assign biasIn_0_w97 = valid0 ? biasIn_0_r30 : wireOut_w97;
assign biasIn_0_w98 = valid0 ? biasIn_0_r29 : wireOut_w98;
assign biasIn_0_w99 = valid0 ? biasIn_0_r28 : wireOut_w99;
assign biasIn_0_w100 = valid0 ? biasIn_0_r27 : wireOut_w100;
assign biasIn_0_w101 = valid0 ? biasIn_0_r26 : wireOut_w101;
assign biasIn_0_w102 = valid0 ? biasIn_0_r25 : wireOut_w102;
assign biasIn_0_w103 = valid0 ? biasIn_0_r24 : wireOut_w103;
assign biasIn_0_w104 = valid0 ? biasIn_0_r23 : wireOut_w104;
assign biasIn_0_w105 = valid0 ? biasIn_0_r22 : wireOut_w105;
assign biasIn_0_w106 = valid0 ? biasIn_0_r21 : wireOut_w106;
assign biasIn_0_w107 = valid0 ? biasIn_0_r20 : wireOut_w107;
assign biasIn_0_w108 = valid0 ? biasIn_0_r19 : wireOut_w108;
assign biasIn_0_w109 = valid0 ? biasIn_0_r18 : wireOut_w109;
assign biasIn_0_w110 = valid0 ? biasIn_0_r17 : wireOut_w110;
assign biasIn_0_w111 = valid0 ? biasIn_0_r16 : wireOut_w111;
assign biasIn_0_w112 = valid0 ? biasIn_0_r15 : wireOut_w112;
assign biasIn_0_w113 = valid0 ? biasIn_0_r14 : wireOut_w113;
assign biasIn_0_w114 = valid0 ? biasIn_0_r13 : wireOut_w114;
assign biasIn_0_w115 = valid0 ? biasIn_0_r12 : wireOut_w115;
assign biasIn_0_w116 = valid0 ? biasIn_0_r11 : wireOut_w116;
assign biasIn_0_w117 = valid0 ? biasIn_0_r10 : wireOut_w117;
assign biasIn_0_w118 = valid0 ? biasIn_0_r9 : wireOut_w118;
assign biasIn_0_w119 = valid0 ? biasIn_0_r8 : wireOut_w119;
assign biasIn_0_w120 = valid0 ? biasIn_0_r7 : wireOut_w120;
assign biasIn_0_w121 = valid0 ? biasIn_0_r6 : wireOut_w121;
assign biasIn_0_w122 = valid0 ? biasIn_0_r5 : wireOut_w122;
assign biasIn_0_w123 = valid0 ? biasIn_0_r4 : wireOut_w123;
assign biasIn_0_w124 = valid0 ? biasIn_0_r3 : wireOut_w124;
assign biasIn_0_w125 = valid0 ? biasIn_0_r2 : wireOut_w125;
assign biasIn_0_w126 = valid0 ? biasIn_0_r1 : wireOut_w126;
assign biasIn_0_w127 = valid0 ? biasIn_0 : wireOut_w127;

// Create the output Delay Line

always @(posedge clk) begin
  if (reset) begin
    outLine_w0 <= 'd0;
    outLine_w1 <= 'd0;
    outLine_w10 <= 'd0;
    outLine_w100 <= 'd0;
    outLine_w101 <= 'd0;
    outLine_w102 <= 'd0;
    outLine_w103 <= 'd0;
    outLine_w104 <= 'd0;
    outLine_w105 <= 'd0;
    outLine_w106 <= 'd0;
    outLine_w107 <= 'd0;
    outLine_w108 <= 'd0;
    outLine_w109 <= 'd0;
    outLine_w11 <= 'd0;
    outLine_w110 <= 'd0;
    outLine_w111 <= 'd0;
    outLine_w112 <= 'd0;
    outLine_w113 <= 'd0;
    outLine_w114 <= 'd0;
    outLine_w115 <= 'd0;
    outLine_w116 <= 'd0;
    outLine_w117 <= 'd0;
    outLine_w118 <= 'd0;
    outLine_w119 <= 'd0;
    outLine_w12 <= 'd0;
    outLine_w120 <= 'd0;
    outLine_w121 <= 'd0;
    outLine_w122 <= 'd0;
    outLine_w123 <= 'd0;
    outLine_w124 <= 'd0;
    outLine_w125 <= 'd0;
    outLine_w126 <= 'd0;
    outLine_w127 <= 'd0;
    outLine_w13 <= 'd0;
    outLine_w14 <= 'd0;
    outLine_w15 <= 'd0;
    outLine_w16 <= 'd0;
    outLine_w17 <= 'd0;
    outLine_w18 <= 'd0;
    outLine_w19 <= 'd0;
    outLine_w2 <= 'd0;
    outLine_w20 <= 'd0;
    outLine_w21 <= 'd0;
    outLine_w22 <= 'd0;
    outLine_w23 <= 'd0;
    outLine_w24 <= 'd0;
    outLine_w25 <= 'd0;
    outLine_w26 <= 'd0;
    outLine_w27 <= 'd0;
    outLine_w28 <= 'd0;
    outLine_w29 <= 'd0;
    outLine_w3 <= 'd0;
    outLine_w30 <= 'd0;
    outLine_w31 <= 'd0;
    outLine_w32 <= 'd0;
    outLine_w33 <= 'd0;
    outLine_w34 <= 'd0;
    outLine_w35 <= 'd0;
    outLine_w36 <= 'd0;
    outLine_w37 <= 'd0;
    outLine_w38 <= 'd0;
    outLine_w39 <= 'd0;
    outLine_w4 <= 'd0;
    outLine_w40 <= 'd0;
    outLine_w41 <= 'd0;
    outLine_w42 <= 'd0;
    outLine_w43 <= 'd0;
    outLine_w44 <= 'd0;
    outLine_w45 <= 'd0;
    outLine_w46 <= 'd0;
    outLine_w47 <= 'd0;
    outLine_w48 <= 'd0;
    outLine_w49 <= 'd0;
    outLine_w5 <= 'd0;
    outLine_w50 <= 'd0;
    outLine_w51 <= 'd0;
    outLine_w52 <= 'd0;
    outLine_w53 <= 'd0;
    outLine_w54 <= 'd0;
    outLine_w55 <= 'd0;
    outLine_w56 <= 'd0;
    outLine_w57 <= 'd0;
    outLine_w58 <= 'd0;
    outLine_w59 <= 'd0;
    outLine_w6 <= 'd0;
    outLine_w60 <= 'd0;
    outLine_w61 <= 'd0;
    outLine_w62 <= 'd0;
    outLine_w63 <= 'd0;
    outLine_w64 <= 'd0;
    outLine_w65 <= 'd0;
    outLine_w66 <= 'd0;
    outLine_w67 <= 'd0;
    outLine_w68 <= 'd0;
    outLine_w69 <= 'd0;
    outLine_w7 <= 'd0;
    outLine_w70 <= 'd0;
    outLine_w71 <= 'd0;
    outLine_w72 <= 'd0;
    outLine_w73 <= 'd0;
    outLine_w74 <= 'd0;
    outLine_w75 <= 'd0;
    outLine_w76 <= 'd0;
    outLine_w77 <= 'd0;
    outLine_w78 <= 'd0;
    outLine_w79 <= 'd0;
    outLine_w8 <= 'd0;
    outLine_w80 <= 'd0;
    outLine_w81 <= 'd0;
    outLine_w82 <= 'd0;
    outLine_w83 <= 'd0;
    outLine_w84 <= 'd0;
    outLine_w85 <= 'd0;
    outLine_w86 <= 'd0;
    outLine_w87 <= 'd0;
    outLine_w88 <= 'd0;
    outLine_w89 <= 'd0;
    outLine_w9 <= 'd0;
    outLine_w90 <= 'd0;
    outLine_w91 <= 'd0;
    outLine_w92 <= 'd0;
    outLine_w93 <= 'd0;
    outLine_w94 <= 'd0;
    outLine_w95 <= 'd0;
    outLine_w96 <= 'd0;
    outLine_w97 <= 'd0;
    outLine_w98 <= 'd0;
    outLine_w99 <= 'd0;
  end
  else begin
    if (valid0) begin
      outLine_w0 <= wireOut_w0;
      outLine_w1 <= wireOut_w1;
      outLine_w2 <= wireOut_w2;
      outLine_w3 <= wireOut_w3;
      outLine_w4 <= wireOut_w4;
      outLine_w5 <= wireOut_w5;
      outLine_w6 <= wireOut_w6;
      outLine_w7 <= wireOut_w7;
      outLine_w8 <= wireOut_w8;
      outLine_w9 <= wireOut_w9;
      outLine_w10 <= wireOut_w10;
      outLine_w11 <= wireOut_w11;
      outLine_w12 <= wireOut_w12;
      outLine_w13 <= wireOut_w13;
      outLine_w14 <= wireOut_w14;
      outLine_w15 <= wireOut_w15;
      outLine_w16 <= wireOut_w16;
      outLine_w17 <= wireOut_w17;
      outLine_w18 <= wireOut_w18;
      outLine_w19 <= wireOut_w19;
      outLine_w20 <= wireOut_w20;
      outLine_w21 <= wireOut_w21;
      outLine_w22 <= wireOut_w22;
      outLine_w23 <= wireOut_w23;
      outLine_w24 <= wireOut_w24;
      outLine_w25 <= wireOut_w25;
      outLine_w26 <= wireOut_w26;
      outLine_w27 <= wireOut_w27;
      outLine_w28 <= wireOut_w28;
      outLine_w29 <= wireOut_w29;
      outLine_w30 <= wireOut_w30;
      outLine_w31 <= wireOut_w31;
      outLine_w32 <= wireOut_w32;
      outLine_w33 <= wireOut_w33;
      outLine_w34 <= wireOut_w34;
      outLine_w35 <= wireOut_w35;
      outLine_w36 <= wireOut_w36;
      outLine_w37 <= wireOut_w37;
      outLine_w38 <= wireOut_w38;
      outLine_w39 <= wireOut_w39;
      outLine_w40 <= wireOut_w40;
      outLine_w41 <= wireOut_w41;
      outLine_w42 <= wireOut_w42;
      outLine_w43 <= wireOut_w43;
      outLine_w44 <= wireOut_w44;
      outLine_w45 <= wireOut_w45;
      outLine_w46 <= wireOut_w46;
      outLine_w47 <= wireOut_w47;
      outLine_w48 <= wireOut_w48;
      outLine_w49 <= wireOut_w49;
      outLine_w50 <= wireOut_w50;
      outLine_w51 <= wireOut_w51;
      outLine_w52 <= wireOut_w52;
      outLine_w53 <= wireOut_w53;
      outLine_w54 <= wireOut_w54;
      outLine_w55 <= wireOut_w55;
      outLine_w56 <= wireOut_w56;
      outLine_w57 <= wireOut_w57;
      outLine_w58 <= wireOut_w58;
      outLine_w59 <= wireOut_w59;
      outLine_w60 <= wireOut_w60;
      outLine_w61 <= wireOut_w61;
      outLine_w62 <= wireOut_w62;
      outLine_w63 <= wireOut_w63;
      outLine_w64 <= wireOut_w64;
      outLine_w65 <= wireOut_w65;
      outLine_w66 <= wireOut_w66;
      outLine_w67 <= wireOut_w67;
      outLine_w68 <= wireOut_w68;
      outLine_w69 <= wireOut_w69;
      outLine_w70 <= wireOut_w70;
      outLine_w71 <= wireOut_w71;
      outLine_w72 <= wireOut_w72;
      outLine_w73 <= wireOut_w73;
      outLine_w74 <= wireOut_w74;
      outLine_w75 <= wireOut_w75;
      outLine_w76 <= wireOut_w76;
      outLine_w77 <= wireOut_w77;
      outLine_w78 <= wireOut_w78;
      outLine_w79 <= wireOut_w79;
      outLine_w80 <= wireOut_w80;
      outLine_w81 <= wireOut_w81;
      outLine_w82 <= wireOut_w82;
      outLine_w83 <= wireOut_w83;
      outLine_w84 <= wireOut_w84;
      outLine_w85 <= wireOut_w85;
      outLine_w86 <= wireOut_w86;
      outLine_w87 <= wireOut_w87;
      outLine_w88 <= wireOut_w88;
      outLine_w89 <= wireOut_w89;
      outLine_w90 <= wireOut_w90;
      outLine_w91 <= wireOut_w91;
      outLine_w92 <= wireOut_w92;
      outLine_w93 <= wireOut_w93;
      outLine_w94 <= wireOut_w94;
      outLine_w95 <= wireOut_w95;
      outLine_w96 <= wireOut_w96;
      outLine_w97 <= wireOut_w97;
      outLine_w98 <= wireOut_w98;
      outLine_w99 <= wireOut_w99;
      outLine_w100 <= wireOut_w100;
      outLine_w101 <= wireOut_w101;
      outLine_w102 <= wireOut_w102;
      outLine_w103 <= wireOut_w103;
      outLine_w104 <= wireOut_w104;
      outLine_w105 <= wireOut_w105;
      outLine_w106 <= wireOut_w106;
      outLine_w107 <= wireOut_w107;
      outLine_w108 <= wireOut_w108;
      outLine_w109 <= wireOut_w109;
      outLine_w110 <= wireOut_w110;
      outLine_w111 <= wireOut_w111;
      outLine_w112 <= wireOut_w112;
      outLine_w113 <= wireOut_w113;
      outLine_w114 <= wireOut_w114;
      outLine_w115 <= wireOut_w115;
      outLine_w116 <= wireOut_w116;
      outLine_w117 <= wireOut_w117;
      outLine_w118 <= wireOut_w118;
      outLine_w119 <= wireOut_w119;
      outLine_w120 <= wireOut_w120;
      outLine_w121 <= wireOut_w121;
      outLine_w122 <= wireOut_w122;
      outLine_w123 <= wireOut_w123;
      outLine_w124 <= wireOut_w124;
      outLine_w125 <= wireOut_w125;
      outLine_w126 <= wireOut_w126;
      outLine_w127 <= wireOut_w127;
    end
    else begin
      outLine_w0 <= outLine_w1;
      outLine_w1 <= outLine_w2;
      outLine_w2 <= outLine_w3;
      outLine_w3 <= outLine_w4;
      outLine_w4 <= outLine_w5;
      outLine_w5 <= outLine_w6;
      outLine_w6 <= outLine_w7;
      outLine_w7 <= outLine_w8;
      outLine_w8 <= outLine_w9;
      outLine_w9 <= outLine_w10;
      outLine_w10 <= outLine_w11;
      outLine_w11 <= outLine_w12;
      outLine_w12 <= outLine_w13;
      outLine_w13 <= outLine_w14;
      outLine_w14 <= outLine_w15;
      outLine_w15 <= outLine_w16;
      outLine_w16 <= outLine_w17;
      outLine_w17 <= outLine_w18;
      outLine_w18 <= outLine_w19;
      outLine_w19 <= outLine_w20;
      outLine_w20 <= outLine_w21;
      outLine_w21 <= outLine_w22;
      outLine_w22 <= outLine_w23;
      outLine_w23 <= outLine_w24;
      outLine_w24 <= outLine_w25;
      outLine_w25 <= outLine_w26;
      outLine_w26 <= outLine_w27;
      outLine_w27 <= outLine_w28;
      outLine_w28 <= outLine_w29;
      outLine_w29 <= outLine_w30;
      outLine_w30 <= outLine_w31;
      outLine_w31 <= outLine_w32;
      outLine_w32 <= outLine_w33;
      outLine_w33 <= outLine_w34;
      outLine_w34 <= outLine_w35;
      outLine_w35 <= outLine_w36;
      outLine_w36 <= outLine_w37;
      outLine_w37 <= outLine_w38;
      outLine_w38 <= outLine_w39;
      outLine_w39 <= outLine_w40;
      outLine_w40 <= outLine_w41;
      outLine_w41 <= outLine_w42;
      outLine_w42 <= outLine_w43;
      outLine_w43 <= outLine_w44;
      outLine_w44 <= outLine_w45;
      outLine_w45 <= outLine_w46;
      outLine_w46 <= outLine_w47;
      outLine_w47 <= outLine_w48;
      outLine_w48 <= outLine_w49;
      outLine_w49 <= outLine_w50;
      outLine_w50 <= outLine_w51;
      outLine_w51 <= outLine_w52;
      outLine_w52 <= outLine_w53;
      outLine_w53 <= outLine_w54;
      outLine_w54 <= outLine_w55;
      outLine_w55 <= outLine_w56;
      outLine_w56 <= outLine_w57;
      outLine_w57 <= outLine_w58;
      outLine_w58 <= outLine_w59;
      outLine_w59 <= outLine_w60;
      outLine_w60 <= outLine_w61;
      outLine_w61 <= outLine_w62;
      outLine_w62 <= outLine_w63;
      outLine_w63 <= outLine_w64;
      outLine_w64 <= outLine_w65;
      outLine_w65 <= outLine_w66;
      outLine_w66 <= outLine_w67;
      outLine_w67 <= outLine_w68;
      outLine_w68 <= outLine_w69;
      outLine_w69 <= outLine_w70;
      outLine_w70 <= outLine_w71;
      outLine_w71 <= outLine_w72;
      outLine_w72 <= outLine_w73;
      outLine_w73 <= outLine_w74;
      outLine_w74 <= outLine_w75;
      outLine_w75 <= outLine_w76;
      outLine_w76 <= outLine_w77;
      outLine_w77 <= outLine_w78;
      outLine_w78 <= outLine_w79;
      outLine_w79 <= outLine_w80;
      outLine_w80 <= outLine_w81;
      outLine_w81 <= outLine_w82;
      outLine_w82 <= outLine_w83;
      outLine_w83 <= outLine_w84;
      outLine_w84 <= outLine_w85;
      outLine_w85 <= outLine_w86;
      outLine_w86 <= outLine_w87;
      outLine_w87 <= outLine_w88;
      outLine_w88 <= outLine_w89;
      outLine_w89 <= outLine_w90;
      outLine_w90 <= outLine_w91;
      outLine_w91 <= outLine_w92;
      outLine_w92 <= outLine_w93;
      outLine_w93 <= outLine_w94;
      outLine_w94 <= outLine_w95;
      outLine_w95 <= outLine_w96;
      outLine_w96 <= outLine_w97;
      outLine_w97 <= outLine_w98;
      outLine_w98 <= outLine_w99;
      outLine_w99 <= outLine_w100;
      outLine_w100 <= outLine_w101;
      outLine_w101 <= outLine_w102;
      outLine_w102 <= outLine_w103;
      outLine_w103 <= outLine_w104;
      outLine_w104 <= outLine_w105;
      outLine_w105 <= outLine_w106;
      outLine_w106 <= outLine_w107;
      outLine_w107 <= outLine_w108;
      outLine_w108 <= outLine_w109;
      outLine_w109 <= outLine_w110;
      outLine_w110 <= outLine_w111;
      outLine_w111 <= outLine_w112;
      outLine_w112 <= outLine_w113;
      outLine_w113 <= outLine_w114;
      outLine_w114 <= outLine_w115;
      outLine_w115 <= outLine_w116;
      outLine_w116 <= outLine_w117;
      outLine_w117 <= outLine_w118;
      outLine_w118 <= outLine_w119;
      outLine_w119 <= outLine_w120;
      outLine_w120 <= outLine_w121;
      outLine_w121 <= outLine_w122;
      outLine_w122 <= outLine_w123;
      outLine_w123 <= outLine_w124;
      outLine_w124 <= outLine_w125;
      outLine_w125 <= outLine_w126;
      outLine_w126 <= outLine_w127;
    end
  end
end

// Assign the outputs
assign dataOutPre_0 = outLine_w0;
endmodule

