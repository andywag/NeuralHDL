//-----------------------------------------------------------------------------
// Company: 			                                                              
// Author:				Andy                                                          
// Date:                                                                       
// Module Name:       testNeuronStage
// Description:                                                                
//                                                                             
//-----------------------------------------------------------------------------
`timescale 10ns/1ns


`ifndef TYPES
  `include "types.v"
  `define TYPES
`endif

    module testNeuronStage(
  input                         clk,
  input                         reset);

// Parameters 



// Wires 

  wire                  [30:0]  d_index           ;  // <31,0>


// Registers 

  reg                   [31:0]  biasIn_0_mem[0:49920];  // <32,0>
  reg                   [31:0]  counter           ;  // <32,0>
  reg                   [31:0]  dataIn_0_mem[0:49920];  // <32,0>
  reg                   [31:0]  rout1_fptr        ;  // <32,0>
  reg                   [31:0]  tapIn_0_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_100_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_101_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_102_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_103_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_104_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_105_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_106_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_107_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_108_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_109_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_10_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_110_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_111_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_112_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_113_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_114_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_115_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_116_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_117_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_118_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_119_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_11_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_120_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_121_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_122_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_123_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_124_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_125_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_126_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_127_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_12_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_13_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_14_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_15_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_16_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_17_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_18_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_19_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_1_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_20_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_21_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_22_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_23_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_24_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_25_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_26_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_27_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_28_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_29_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_2_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_30_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_31_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_32_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_33_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_34_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_35_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_36_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_37_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_38_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_39_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_3_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_40_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_41_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_42_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_43_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_44_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_45_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_46_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_47_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_48_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_49_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_4_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_50_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_51_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_52_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_53_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_54_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_55_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_56_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_57_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_58_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_59_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_5_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_60_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_61_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_62_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_63_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_64_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_65_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_66_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_67_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_68_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_69_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_6_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_70_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_71_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_72_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_73_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_74_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_75_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_76_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_77_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_78_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_79_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_7_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_80_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_81_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_82_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_83_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_84_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_85_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_86_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_87_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_88_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_89_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_8_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_90_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_91_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_92_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_93_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_94_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_95_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_96_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_97_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_98_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_99_mem[0:6389760];  // <32,0>
  reg                   [31:0]  tapIn_9_mem[0:6389760];  // <32,0>
  reg                           valid             ;  // <1,0>


// Other

  float_24_8                    biasIn_0;  // <1,0>
  float_24_8                    biasIn_0_0;  // <1,0>
  float_24_8                    biasIn_0_1;  // <1,0>
  float_24_8                    biasIn_0_10;  // <1,0>
  float_24_8                    biasIn_0_100;  // <1,0>
  float_24_8                    biasIn_0_101;  // <1,0>
  float_24_8                    biasIn_0_102;  // <1,0>
  float_24_8                    biasIn_0_103;  // <1,0>
  float_24_8                    biasIn_0_104;  // <1,0>
  float_24_8                    biasIn_0_105;  // <1,0>
  float_24_8                    biasIn_0_106;  // <1,0>
  float_24_8                    biasIn_0_107;  // <1,0>
  float_24_8                    biasIn_0_108;  // <1,0>
  float_24_8                    biasIn_0_109;  // <1,0>
  float_24_8                    biasIn_0_11;  // <1,0>
  float_24_8                    biasIn_0_110;  // <1,0>
  float_24_8                    biasIn_0_111;  // <1,0>
  float_24_8                    biasIn_0_112;  // <1,0>
  float_24_8                    biasIn_0_113;  // <1,0>
  float_24_8                    biasIn_0_114;  // <1,0>
  float_24_8                    biasIn_0_115;  // <1,0>
  float_24_8                    biasIn_0_116;  // <1,0>
  float_24_8                    biasIn_0_117;  // <1,0>
  float_24_8                    biasIn_0_118;  // <1,0>
  float_24_8                    biasIn_0_119;  // <1,0>
  float_24_8                    biasIn_0_12;  // <1,0>
  float_24_8                    biasIn_0_120;  // <1,0>
  float_24_8                    biasIn_0_121;  // <1,0>
  float_24_8                    biasIn_0_122;  // <1,0>
  float_24_8                    biasIn_0_123;  // <1,0>
  float_24_8                    biasIn_0_124;  // <1,0>
  float_24_8                    biasIn_0_125;  // <1,0>
  float_24_8                    biasIn_0_126;  // <1,0>
  float_24_8                    biasIn_0_127;  // <1,0>
  float_24_8                    biasIn_0_13;  // <1,0>
  float_24_8                    biasIn_0_14;  // <1,0>
  float_24_8                    biasIn_0_15;  // <1,0>
  float_24_8                    biasIn_0_16;  // <1,0>
  float_24_8                    biasIn_0_17;  // <1,0>
  float_24_8                    biasIn_0_18;  // <1,0>
  float_24_8                    biasIn_0_19;  // <1,0>
  float_24_8                    biasIn_0_2;  // <1,0>
  float_24_8                    biasIn_0_20;  // <1,0>
  float_24_8                    biasIn_0_21;  // <1,0>
  float_24_8                    biasIn_0_22;  // <1,0>
  float_24_8                    biasIn_0_23;  // <1,0>
  float_24_8                    biasIn_0_24;  // <1,0>
  float_24_8                    biasIn_0_25;  // <1,0>
  float_24_8                    biasIn_0_26;  // <1,0>
  float_24_8                    biasIn_0_27;  // <1,0>
  float_24_8                    biasIn_0_28;  // <1,0>
  float_24_8                    biasIn_0_29;  // <1,0>
  float_24_8                    biasIn_0_3;  // <1,0>
  float_24_8                    biasIn_0_30;  // <1,0>
  float_24_8                    biasIn_0_31;  // <1,0>
  float_24_8                    biasIn_0_32;  // <1,0>
  float_24_8                    biasIn_0_33;  // <1,0>
  float_24_8                    biasIn_0_34;  // <1,0>
  float_24_8                    biasIn_0_35;  // <1,0>
  float_24_8                    biasIn_0_36;  // <1,0>
  float_24_8                    biasIn_0_37;  // <1,0>
  float_24_8                    biasIn_0_38;  // <1,0>
  float_24_8                    biasIn_0_39;  // <1,0>
  float_24_8                    biasIn_0_4;  // <1,0>
  float_24_8                    biasIn_0_40;  // <1,0>
  float_24_8                    biasIn_0_41;  // <1,0>
  float_24_8                    biasIn_0_42;  // <1,0>
  float_24_8                    biasIn_0_43;  // <1,0>
  float_24_8                    biasIn_0_44;  // <1,0>
  float_24_8                    biasIn_0_45;  // <1,0>
  float_24_8                    biasIn_0_46;  // <1,0>
  float_24_8                    biasIn_0_47;  // <1,0>
  float_24_8                    biasIn_0_48;  // <1,0>
  float_24_8                    biasIn_0_49;  // <1,0>
  float_24_8                    biasIn_0_5;  // <1,0>
  float_24_8                    biasIn_0_50;  // <1,0>
  float_24_8                    biasIn_0_51;  // <1,0>
  float_24_8                    biasIn_0_52;  // <1,0>
  float_24_8                    biasIn_0_53;  // <1,0>
  float_24_8                    biasIn_0_54;  // <1,0>
  float_24_8                    biasIn_0_55;  // <1,0>
  float_24_8                    biasIn_0_56;  // <1,0>
  float_24_8                    biasIn_0_57;  // <1,0>
  float_24_8                    biasIn_0_58;  // <1,0>
  float_24_8                    biasIn_0_59;  // <1,0>
  float_24_8                    biasIn_0_6;  // <1,0>
  float_24_8                    biasIn_0_60;  // <1,0>
  float_24_8                    biasIn_0_61;  // <1,0>
  float_24_8                    biasIn_0_62;  // <1,0>
  float_24_8                    biasIn_0_63;  // <1,0>
  float_24_8                    biasIn_0_64;  // <1,0>
  float_24_8                    biasIn_0_65;  // <1,0>
  float_24_8                    biasIn_0_66;  // <1,0>
  float_24_8                    biasIn_0_67;  // <1,0>
  float_24_8                    biasIn_0_68;  // <1,0>
  float_24_8                    biasIn_0_69;  // <1,0>
  float_24_8                    biasIn_0_7;  // <1,0>
  float_24_8                    biasIn_0_70;  // <1,0>
  float_24_8                    biasIn_0_71;  // <1,0>
  float_24_8                    biasIn_0_72;  // <1,0>
  float_24_8                    biasIn_0_73;  // <1,0>
  float_24_8                    biasIn_0_74;  // <1,0>
  float_24_8                    biasIn_0_75;  // <1,0>
  float_24_8                    biasIn_0_76;  // <1,0>
  float_24_8                    biasIn_0_77;  // <1,0>
  float_24_8                    biasIn_0_78;  // <1,0>
  float_24_8                    biasIn_0_79;  // <1,0>
  float_24_8                    biasIn_0_8;  // <1,0>
  float_24_8                    biasIn_0_80;  // <1,0>
  float_24_8                    biasIn_0_81;  // <1,0>
  float_24_8                    biasIn_0_82;  // <1,0>
  float_24_8                    biasIn_0_83;  // <1,0>
  float_24_8                    biasIn_0_84;  // <1,0>
  float_24_8                    biasIn_0_85;  // <1,0>
  float_24_8                    biasIn_0_86;  // <1,0>
  float_24_8                    biasIn_0_87;  // <1,0>
  float_24_8                    biasIn_0_88;  // <1,0>
  float_24_8                    biasIn_0_89;  // <1,0>
  float_24_8                    biasIn_0_9;  // <1,0>
  float_24_8                    biasIn_0_90;  // <1,0>
  float_24_8                    biasIn_0_91;  // <1,0>
  float_24_8                    biasIn_0_92;  // <1,0>
  float_24_8                    biasIn_0_93;  // <1,0>
  float_24_8                    biasIn_0_94;  // <1,0>
  float_24_8                    biasIn_0_95;  // <1,0>
  float_24_8                    biasIn_0_96;  // <1,0>
  float_24_8                    biasIn_0_97;  // <1,0>
  float_24_8                    biasIn_0_98;  // <1,0>
  float_24_8                    biasIn_0_99;  // <1,0>
  float_24_8                    dataIn_0;  // <1,0>
  float_24_8                    dataOutPre_0;  // <1,0>
  float_24_8                    dataOut_0;  // <1,0>
  float_24_8                    tapIn_0;  // <1,0>
  float_24_8                    tapIn_1;  // <1,0>
  float_24_8                    tapIn_10;  // <1,0>
  float_24_8                    tapIn_100;  // <1,0>
  float_24_8                    tapIn_101;  // <1,0>
  float_24_8                    tapIn_102;  // <1,0>
  float_24_8                    tapIn_103;  // <1,0>
  float_24_8                    tapIn_104;  // <1,0>
  float_24_8                    tapIn_105;  // <1,0>
  float_24_8                    tapIn_106;  // <1,0>
  float_24_8                    tapIn_107;  // <1,0>
  float_24_8                    tapIn_108;  // <1,0>
  float_24_8                    tapIn_109;  // <1,0>
  float_24_8                    tapIn_11;  // <1,0>
  float_24_8                    tapIn_110;  // <1,0>
  float_24_8                    tapIn_111;  // <1,0>
  float_24_8                    tapIn_112;  // <1,0>
  float_24_8                    tapIn_113;  // <1,0>
  float_24_8                    tapIn_114;  // <1,0>
  float_24_8                    tapIn_115;  // <1,0>
  float_24_8                    tapIn_116;  // <1,0>
  float_24_8                    tapIn_117;  // <1,0>
  float_24_8                    tapIn_118;  // <1,0>
  float_24_8                    tapIn_119;  // <1,0>
  float_24_8                    tapIn_12;  // <1,0>
  float_24_8                    tapIn_120;  // <1,0>
  float_24_8                    tapIn_121;  // <1,0>
  float_24_8                    tapIn_122;  // <1,0>
  float_24_8                    tapIn_123;  // <1,0>
  float_24_8                    tapIn_124;  // <1,0>
  float_24_8                    tapIn_125;  // <1,0>
  float_24_8                    tapIn_126;  // <1,0>
  float_24_8                    tapIn_127;  // <1,0>
  float_24_8                    tapIn_13;  // <1,0>
  float_24_8                    tapIn_14;  // <1,0>
  float_24_8                    tapIn_15;  // <1,0>
  float_24_8                    tapIn_16;  // <1,0>
  float_24_8                    tapIn_17;  // <1,0>
  float_24_8                    tapIn_18;  // <1,0>
  float_24_8                    tapIn_19;  // <1,0>
  float_24_8                    tapIn_2;  // <1,0>
  float_24_8                    tapIn_20;  // <1,0>
  float_24_8                    tapIn_21;  // <1,0>
  float_24_8                    tapIn_22;  // <1,0>
  float_24_8                    tapIn_23;  // <1,0>
  float_24_8                    tapIn_24;  // <1,0>
  float_24_8                    tapIn_25;  // <1,0>
  float_24_8                    tapIn_26;  // <1,0>
  float_24_8                    tapIn_27;  // <1,0>
  float_24_8                    tapIn_28;  // <1,0>
  float_24_8                    tapIn_29;  // <1,0>
  float_24_8                    tapIn_3;  // <1,0>
  float_24_8                    tapIn_30;  // <1,0>
  float_24_8                    tapIn_31;  // <1,0>
  float_24_8                    tapIn_32;  // <1,0>
  float_24_8                    tapIn_33;  // <1,0>
  float_24_8                    tapIn_34;  // <1,0>
  float_24_8                    tapIn_35;  // <1,0>
  float_24_8                    tapIn_36;  // <1,0>
  float_24_8                    tapIn_37;  // <1,0>
  float_24_8                    tapIn_38;  // <1,0>
  float_24_8                    tapIn_39;  // <1,0>
  float_24_8                    tapIn_4;  // <1,0>
  float_24_8                    tapIn_40;  // <1,0>
  float_24_8                    tapIn_41;  // <1,0>
  float_24_8                    tapIn_42;  // <1,0>
  float_24_8                    tapIn_43;  // <1,0>
  float_24_8                    tapIn_44;  // <1,0>
  float_24_8                    tapIn_45;  // <1,0>
  float_24_8                    tapIn_46;  // <1,0>
  float_24_8                    tapIn_47;  // <1,0>
  float_24_8                    tapIn_48;  // <1,0>
  float_24_8                    tapIn_49;  // <1,0>
  float_24_8                    tapIn_5;  // <1,0>
  float_24_8                    tapIn_50;  // <1,0>
  float_24_8                    tapIn_51;  // <1,0>
  float_24_8                    tapIn_52;  // <1,0>
  float_24_8                    tapIn_53;  // <1,0>
  float_24_8                    tapIn_54;  // <1,0>
  float_24_8                    tapIn_55;  // <1,0>
  float_24_8                    tapIn_56;  // <1,0>
  float_24_8                    tapIn_57;  // <1,0>
  float_24_8                    tapIn_58;  // <1,0>
  float_24_8                    tapIn_59;  // <1,0>
  float_24_8                    tapIn_6;  // <1,0>
  float_24_8                    tapIn_60;  // <1,0>
  float_24_8                    tapIn_61;  // <1,0>
  float_24_8                    tapIn_62;  // <1,0>
  float_24_8                    tapIn_63;  // <1,0>
  float_24_8                    tapIn_64;  // <1,0>
  float_24_8                    tapIn_65;  // <1,0>
  float_24_8                    tapIn_66;  // <1,0>
  float_24_8                    tapIn_67;  // <1,0>
  float_24_8                    tapIn_68;  // <1,0>
  float_24_8                    tapIn_69;  // <1,0>
  float_24_8                    tapIn_7;  // <1,0>
  float_24_8                    tapIn_70;  // <1,0>
  float_24_8                    tapIn_71;  // <1,0>
  float_24_8                    tapIn_72;  // <1,0>
  float_24_8                    tapIn_73;  // <1,0>
  float_24_8                    tapIn_74;  // <1,0>
  float_24_8                    tapIn_75;  // <1,0>
  float_24_8                    tapIn_76;  // <1,0>
  float_24_8                    tapIn_77;  // <1,0>
  float_24_8                    tapIn_78;  // <1,0>
  float_24_8                    tapIn_79;  // <1,0>
  float_24_8                    tapIn_8;  // <1,0>
  float_24_8                    tapIn_80;  // <1,0>
  float_24_8                    tapIn_81;  // <1,0>
  float_24_8                    tapIn_82;  // <1,0>
  float_24_8                    tapIn_83;  // <1,0>
  float_24_8                    tapIn_84;  // <1,0>
  float_24_8                    tapIn_85;  // <1,0>
  float_24_8                    tapIn_86;  // <1,0>
  float_24_8                    tapIn_87;  // <1,0>
  float_24_8                    tapIn_88;  // <1,0>
  float_24_8                    tapIn_89;  // <1,0>
  float_24_8                    tapIn_9;  // <1,0>
  float_24_8                    tapIn_90;  // <1,0>
  float_24_8                    tapIn_91;  // <1,0>
  float_24_8                    tapIn_92;  // <1,0>
  float_24_8                    tapIn_93;  // <1,0>
  float_24_8                    tapIn_94;  // <1,0>
  float_24_8                    tapIn_95;  // <1,0>
  float_24_8                    tapIn_96;  // <1,0>
  float_24_8                    tapIn_97;  // <1,0>
  float_24_8                    tapIn_98;  // <1,0>
  float_24_8                    tapIn_99;  // <1,0>


////////////////////////////////////////////////////////////////////////////////
// neuronStage
////////////////////////////////////////////////////////////////////////////////

neuronStage neuronStage (
    .biasIn_0(biasIn_0),
    .clk(clk),
    .dataIn_0(dataIn_0),
    .dataOutPre_0(dataOutPre_0),
    .dataOut_0(dataOut_0),
    .reset(reset),
    .tapIn_0(tapIn_0),
    .tapIn_1(tapIn_1),
    .tapIn_10(tapIn_10),
    .tapIn_100(tapIn_100),
    .tapIn_101(tapIn_101),
    .tapIn_102(tapIn_102),
    .tapIn_103(tapIn_103),
    .tapIn_104(tapIn_104),
    .tapIn_105(tapIn_105),
    .tapIn_106(tapIn_106),
    .tapIn_107(tapIn_107),
    .tapIn_108(tapIn_108),
    .tapIn_109(tapIn_109),
    .tapIn_11(tapIn_11),
    .tapIn_110(tapIn_110),
    .tapIn_111(tapIn_111),
    .tapIn_112(tapIn_112),
    .tapIn_113(tapIn_113),
    .tapIn_114(tapIn_114),
    .tapIn_115(tapIn_115),
    .tapIn_116(tapIn_116),
    .tapIn_117(tapIn_117),
    .tapIn_118(tapIn_118),
    .tapIn_119(tapIn_119),
    .tapIn_12(tapIn_12),
    .tapIn_120(tapIn_120),
    .tapIn_121(tapIn_121),
    .tapIn_122(tapIn_122),
    .tapIn_123(tapIn_123),
    .tapIn_124(tapIn_124),
    .tapIn_125(tapIn_125),
    .tapIn_126(tapIn_126),
    .tapIn_127(tapIn_127),
    .tapIn_13(tapIn_13),
    .tapIn_14(tapIn_14),
    .tapIn_15(tapIn_15),
    .tapIn_16(tapIn_16),
    .tapIn_17(tapIn_17),
    .tapIn_18(tapIn_18),
    .tapIn_19(tapIn_19),
    .tapIn_2(tapIn_2),
    .tapIn_20(tapIn_20),
    .tapIn_21(tapIn_21),
    .tapIn_22(tapIn_22),
    .tapIn_23(tapIn_23),
    .tapIn_24(tapIn_24),
    .tapIn_25(tapIn_25),
    .tapIn_26(tapIn_26),
    .tapIn_27(tapIn_27),
    .tapIn_28(tapIn_28),
    .tapIn_29(tapIn_29),
    .tapIn_3(tapIn_3),
    .tapIn_30(tapIn_30),
    .tapIn_31(tapIn_31),
    .tapIn_32(tapIn_32),
    .tapIn_33(tapIn_33),
    .tapIn_34(tapIn_34),
    .tapIn_35(tapIn_35),
    .tapIn_36(tapIn_36),
    .tapIn_37(tapIn_37),
    .tapIn_38(tapIn_38),
    .tapIn_39(tapIn_39),
    .tapIn_4(tapIn_4),
    .tapIn_40(tapIn_40),
    .tapIn_41(tapIn_41),
    .tapIn_42(tapIn_42),
    .tapIn_43(tapIn_43),
    .tapIn_44(tapIn_44),
    .tapIn_45(tapIn_45),
    .tapIn_46(tapIn_46),
    .tapIn_47(tapIn_47),
    .tapIn_48(tapIn_48),
    .tapIn_49(tapIn_49),
    .tapIn_5(tapIn_5),
    .tapIn_50(tapIn_50),
    .tapIn_51(tapIn_51),
    .tapIn_52(tapIn_52),
    .tapIn_53(tapIn_53),
    .tapIn_54(tapIn_54),
    .tapIn_55(tapIn_55),
    .tapIn_56(tapIn_56),
    .tapIn_57(tapIn_57),
    .tapIn_58(tapIn_58),
    .tapIn_59(tapIn_59),
    .tapIn_6(tapIn_6),
    .tapIn_60(tapIn_60),
    .tapIn_61(tapIn_61),
    .tapIn_62(tapIn_62),
    .tapIn_63(tapIn_63),
    .tapIn_64(tapIn_64),
    .tapIn_65(tapIn_65),
    .tapIn_66(tapIn_66),
    .tapIn_67(tapIn_67),
    .tapIn_68(tapIn_68),
    .tapIn_69(tapIn_69),
    .tapIn_7(tapIn_7),
    .tapIn_70(tapIn_70),
    .tapIn_71(tapIn_71),
    .tapIn_72(tapIn_72),
    .tapIn_73(tapIn_73),
    .tapIn_74(tapIn_74),
    .tapIn_75(tapIn_75),
    .tapIn_76(tapIn_76),
    .tapIn_77(tapIn_77),
    .tapIn_78(tapIn_78),
    .tapIn_79(tapIn_79),
    .tapIn_8(tapIn_8),
    .tapIn_80(tapIn_80),
    .tapIn_81(tapIn_81),
    .tapIn_82(tapIn_82),
    .tapIn_83(tapIn_83),
    .tapIn_84(tapIn_84),
    .tapIn_85(tapIn_85),
    .tapIn_86(tapIn_86),
    .tapIn_87(tapIn_87),
    .tapIn_88(tapIn_88),
    .tapIn_89(tapIn_89),
    .tapIn_9(tapIn_9),
    .tapIn_90(tapIn_90),
    .tapIn_91(tapIn_91),
    .tapIn_92(tapIn_92),
    .tapIn_93(tapIn_93),
    .tapIn_94(tapIn_94),
    .tapIn_95(tapIn_95),
    .tapIn_96(tapIn_96),
    .tapIn_97(tapIn_97),
    .tapIn_98(tapIn_98),
    .tapIn_99(tapIn_99),
    .valid(valid));


// Stop the test when the data runs out
always @(posedge clk) begin
  if (reset) begin
    
  end
  else begin
    if ((counter == 'd50000)) begin
      $finish;
    end
  end
end

// Create a valid pulse
assign valid = (counter[6:0] == 'd126);

// Delay the bias to line up the data
assign d_index = counter[30:0] - 31'd126;

// Load dataIn_0
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/data.hex",dataIn_0_mem);
end

assign dataIn_0 = dataIn_0_mem[d_index];

// Load tapIn_0
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap0.hex",tapIn_0_mem);
end

assign tapIn_0 = tapIn_0_mem[d_index];

// Load tapIn_1
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap1.hex",tapIn_1_mem);
end

assign tapIn_1 = tapIn_1_mem[d_index];

// Load tapIn_2
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap2.hex",tapIn_2_mem);
end

assign tapIn_2 = tapIn_2_mem[d_index];

// Load tapIn_3
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap3.hex",tapIn_3_mem);
end

assign tapIn_3 = tapIn_3_mem[d_index];

// Load tapIn_4
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap4.hex",tapIn_4_mem);
end

assign tapIn_4 = tapIn_4_mem[d_index];

// Load tapIn_5
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap5.hex",tapIn_5_mem);
end

assign tapIn_5 = tapIn_5_mem[d_index];

// Load tapIn_6
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap6.hex",tapIn_6_mem);
end

assign tapIn_6 = tapIn_6_mem[d_index];

// Load tapIn_7
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap7.hex",tapIn_7_mem);
end

assign tapIn_7 = tapIn_7_mem[d_index];

// Load tapIn_8
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap8.hex",tapIn_8_mem);
end

assign tapIn_8 = tapIn_8_mem[d_index];

// Load tapIn_9
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap9.hex",tapIn_9_mem);
end

assign tapIn_9 = tapIn_9_mem[d_index];

// Load tapIn_10
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap10.hex",tapIn_10_mem);
end

assign tapIn_10 = tapIn_10_mem[d_index];

// Load tapIn_11
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap11.hex",tapIn_11_mem);
end

assign tapIn_11 = tapIn_11_mem[d_index];

// Load tapIn_12
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap12.hex",tapIn_12_mem);
end

assign tapIn_12 = tapIn_12_mem[d_index];

// Load tapIn_13
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap13.hex",tapIn_13_mem);
end

assign tapIn_13 = tapIn_13_mem[d_index];

// Load tapIn_14
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap14.hex",tapIn_14_mem);
end

assign tapIn_14 = tapIn_14_mem[d_index];

// Load tapIn_15
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap15.hex",tapIn_15_mem);
end

assign tapIn_15 = tapIn_15_mem[d_index];

// Load tapIn_16
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap16.hex",tapIn_16_mem);
end

assign tapIn_16 = tapIn_16_mem[d_index];

// Load tapIn_17
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap17.hex",tapIn_17_mem);
end

assign tapIn_17 = tapIn_17_mem[d_index];

// Load tapIn_18
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap18.hex",tapIn_18_mem);
end

assign tapIn_18 = tapIn_18_mem[d_index];

// Load tapIn_19
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap19.hex",tapIn_19_mem);
end

assign tapIn_19 = tapIn_19_mem[d_index];

// Load tapIn_20
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap20.hex",tapIn_20_mem);
end

assign tapIn_20 = tapIn_20_mem[d_index];

// Load tapIn_21
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap21.hex",tapIn_21_mem);
end

assign tapIn_21 = tapIn_21_mem[d_index];

// Load tapIn_22
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap22.hex",tapIn_22_mem);
end

assign tapIn_22 = tapIn_22_mem[d_index];

// Load tapIn_23
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap23.hex",tapIn_23_mem);
end

assign tapIn_23 = tapIn_23_mem[d_index];

// Load tapIn_24
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap24.hex",tapIn_24_mem);
end

assign tapIn_24 = tapIn_24_mem[d_index];

// Load tapIn_25
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap25.hex",tapIn_25_mem);
end

assign tapIn_25 = tapIn_25_mem[d_index];

// Load tapIn_26
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap26.hex",tapIn_26_mem);
end

assign tapIn_26 = tapIn_26_mem[d_index];

// Load tapIn_27
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap27.hex",tapIn_27_mem);
end

assign tapIn_27 = tapIn_27_mem[d_index];

// Load tapIn_28
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap28.hex",tapIn_28_mem);
end

assign tapIn_28 = tapIn_28_mem[d_index];

// Load tapIn_29
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap29.hex",tapIn_29_mem);
end

assign tapIn_29 = tapIn_29_mem[d_index];

// Load tapIn_30
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap30.hex",tapIn_30_mem);
end

assign tapIn_30 = tapIn_30_mem[d_index];

// Load tapIn_31
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap31.hex",tapIn_31_mem);
end

assign tapIn_31 = tapIn_31_mem[d_index];

// Load tapIn_32
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap32.hex",tapIn_32_mem);
end

assign tapIn_32 = tapIn_32_mem[d_index];

// Load tapIn_33
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap33.hex",tapIn_33_mem);
end

assign tapIn_33 = tapIn_33_mem[d_index];

// Load tapIn_34
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap34.hex",tapIn_34_mem);
end

assign tapIn_34 = tapIn_34_mem[d_index];

// Load tapIn_35
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap35.hex",tapIn_35_mem);
end

assign tapIn_35 = tapIn_35_mem[d_index];

// Load tapIn_36
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap36.hex",tapIn_36_mem);
end

assign tapIn_36 = tapIn_36_mem[d_index];

// Load tapIn_37
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap37.hex",tapIn_37_mem);
end

assign tapIn_37 = tapIn_37_mem[d_index];

// Load tapIn_38
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap38.hex",tapIn_38_mem);
end

assign tapIn_38 = tapIn_38_mem[d_index];

// Load tapIn_39
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap39.hex",tapIn_39_mem);
end

assign tapIn_39 = tapIn_39_mem[d_index];

// Load tapIn_40
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap40.hex",tapIn_40_mem);
end

assign tapIn_40 = tapIn_40_mem[d_index];

// Load tapIn_41
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap41.hex",tapIn_41_mem);
end

assign tapIn_41 = tapIn_41_mem[d_index];

// Load tapIn_42
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap42.hex",tapIn_42_mem);
end

assign tapIn_42 = tapIn_42_mem[d_index];

// Load tapIn_43
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap43.hex",tapIn_43_mem);
end

assign tapIn_43 = tapIn_43_mem[d_index];

// Load tapIn_44
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap44.hex",tapIn_44_mem);
end

assign tapIn_44 = tapIn_44_mem[d_index];

// Load tapIn_45
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap45.hex",tapIn_45_mem);
end

assign tapIn_45 = tapIn_45_mem[d_index];

// Load tapIn_46
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap46.hex",tapIn_46_mem);
end

assign tapIn_46 = tapIn_46_mem[d_index];

// Load tapIn_47
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap47.hex",tapIn_47_mem);
end

assign tapIn_47 = tapIn_47_mem[d_index];

// Load tapIn_48
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap48.hex",tapIn_48_mem);
end

assign tapIn_48 = tapIn_48_mem[d_index];

// Load tapIn_49
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap49.hex",tapIn_49_mem);
end

assign tapIn_49 = tapIn_49_mem[d_index];

// Load tapIn_50
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap50.hex",tapIn_50_mem);
end

assign tapIn_50 = tapIn_50_mem[d_index];

// Load tapIn_51
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap51.hex",tapIn_51_mem);
end

assign tapIn_51 = tapIn_51_mem[d_index];

// Load tapIn_52
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap52.hex",tapIn_52_mem);
end

assign tapIn_52 = tapIn_52_mem[d_index];

// Load tapIn_53
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap53.hex",tapIn_53_mem);
end

assign tapIn_53 = tapIn_53_mem[d_index];

// Load tapIn_54
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap54.hex",tapIn_54_mem);
end

assign tapIn_54 = tapIn_54_mem[d_index];

// Load tapIn_55
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap55.hex",tapIn_55_mem);
end

assign tapIn_55 = tapIn_55_mem[d_index];

// Load tapIn_56
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap56.hex",tapIn_56_mem);
end

assign tapIn_56 = tapIn_56_mem[d_index];

// Load tapIn_57
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap57.hex",tapIn_57_mem);
end

assign tapIn_57 = tapIn_57_mem[d_index];

// Load tapIn_58
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap58.hex",tapIn_58_mem);
end

assign tapIn_58 = tapIn_58_mem[d_index];

// Load tapIn_59
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap59.hex",tapIn_59_mem);
end

assign tapIn_59 = tapIn_59_mem[d_index];

// Load tapIn_60
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap60.hex",tapIn_60_mem);
end

assign tapIn_60 = tapIn_60_mem[d_index];

// Load tapIn_61
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap61.hex",tapIn_61_mem);
end

assign tapIn_61 = tapIn_61_mem[d_index];

// Load tapIn_62
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap62.hex",tapIn_62_mem);
end

assign tapIn_62 = tapIn_62_mem[d_index];

// Load tapIn_63
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap63.hex",tapIn_63_mem);
end

assign tapIn_63 = tapIn_63_mem[d_index];

// Load tapIn_64
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap64.hex",tapIn_64_mem);
end

assign tapIn_64 = tapIn_64_mem[d_index];

// Load tapIn_65
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap65.hex",tapIn_65_mem);
end

assign tapIn_65 = tapIn_65_mem[d_index];

// Load tapIn_66
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap66.hex",tapIn_66_mem);
end

assign tapIn_66 = tapIn_66_mem[d_index];

// Load tapIn_67
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap67.hex",tapIn_67_mem);
end

assign tapIn_67 = tapIn_67_mem[d_index];

// Load tapIn_68
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap68.hex",tapIn_68_mem);
end

assign tapIn_68 = tapIn_68_mem[d_index];

// Load tapIn_69
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap69.hex",tapIn_69_mem);
end

assign tapIn_69 = tapIn_69_mem[d_index];

// Load tapIn_70
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap70.hex",tapIn_70_mem);
end

assign tapIn_70 = tapIn_70_mem[d_index];

// Load tapIn_71
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap71.hex",tapIn_71_mem);
end

assign tapIn_71 = tapIn_71_mem[d_index];

// Load tapIn_72
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap72.hex",tapIn_72_mem);
end

assign tapIn_72 = tapIn_72_mem[d_index];

// Load tapIn_73
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap73.hex",tapIn_73_mem);
end

assign tapIn_73 = tapIn_73_mem[d_index];

// Load tapIn_74
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap74.hex",tapIn_74_mem);
end

assign tapIn_74 = tapIn_74_mem[d_index];

// Load tapIn_75
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap75.hex",tapIn_75_mem);
end

assign tapIn_75 = tapIn_75_mem[d_index];

// Load tapIn_76
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap76.hex",tapIn_76_mem);
end

assign tapIn_76 = tapIn_76_mem[d_index];

// Load tapIn_77
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap77.hex",tapIn_77_mem);
end

assign tapIn_77 = tapIn_77_mem[d_index];

// Load tapIn_78
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap78.hex",tapIn_78_mem);
end

assign tapIn_78 = tapIn_78_mem[d_index];

// Load tapIn_79
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap79.hex",tapIn_79_mem);
end

assign tapIn_79 = tapIn_79_mem[d_index];

// Load tapIn_80
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap80.hex",tapIn_80_mem);
end

assign tapIn_80 = tapIn_80_mem[d_index];

// Load tapIn_81
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap81.hex",tapIn_81_mem);
end

assign tapIn_81 = tapIn_81_mem[d_index];

// Load tapIn_82
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap82.hex",tapIn_82_mem);
end

assign tapIn_82 = tapIn_82_mem[d_index];

// Load tapIn_83
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap83.hex",tapIn_83_mem);
end

assign tapIn_83 = tapIn_83_mem[d_index];

// Load tapIn_84
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap84.hex",tapIn_84_mem);
end

assign tapIn_84 = tapIn_84_mem[d_index];

// Load tapIn_85
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap85.hex",tapIn_85_mem);
end

assign tapIn_85 = tapIn_85_mem[d_index];

// Load tapIn_86
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap86.hex",tapIn_86_mem);
end

assign tapIn_86 = tapIn_86_mem[d_index];

// Load tapIn_87
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap87.hex",tapIn_87_mem);
end

assign tapIn_87 = tapIn_87_mem[d_index];

// Load tapIn_88
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap88.hex",tapIn_88_mem);
end

assign tapIn_88 = tapIn_88_mem[d_index];

// Load tapIn_89
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap89.hex",tapIn_89_mem);
end

assign tapIn_89 = tapIn_89_mem[d_index];

// Load tapIn_90
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap90.hex",tapIn_90_mem);
end

assign tapIn_90 = tapIn_90_mem[d_index];

// Load tapIn_91
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap91.hex",tapIn_91_mem);
end

assign tapIn_91 = tapIn_91_mem[d_index];

// Load tapIn_92
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap92.hex",tapIn_92_mem);
end

assign tapIn_92 = tapIn_92_mem[d_index];

// Load tapIn_93
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap93.hex",tapIn_93_mem);
end

assign tapIn_93 = tapIn_93_mem[d_index];

// Load tapIn_94
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap94.hex",tapIn_94_mem);
end

assign tapIn_94 = tapIn_94_mem[d_index];

// Load tapIn_95
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap95.hex",tapIn_95_mem);
end

assign tapIn_95 = tapIn_95_mem[d_index];

// Load tapIn_96
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap96.hex",tapIn_96_mem);
end

assign tapIn_96 = tapIn_96_mem[d_index];

// Load tapIn_97
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap97.hex",tapIn_97_mem);
end

assign tapIn_97 = tapIn_97_mem[d_index];

// Load tapIn_98
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap98.hex",tapIn_98_mem);
end

assign tapIn_98 = tapIn_98_mem[d_index];

// Load tapIn_99
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap99.hex",tapIn_99_mem);
end

assign tapIn_99 = tapIn_99_mem[d_index];

// Load tapIn_100
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap100.hex",tapIn_100_mem);
end

assign tapIn_100 = tapIn_100_mem[d_index];

// Load tapIn_101
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap101.hex",tapIn_101_mem);
end

assign tapIn_101 = tapIn_101_mem[d_index];

// Load tapIn_102
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap102.hex",tapIn_102_mem);
end

assign tapIn_102 = tapIn_102_mem[d_index];

// Load tapIn_103
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap103.hex",tapIn_103_mem);
end

assign tapIn_103 = tapIn_103_mem[d_index];

// Load tapIn_104
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap104.hex",tapIn_104_mem);
end

assign tapIn_104 = tapIn_104_mem[d_index];

// Load tapIn_105
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap105.hex",tapIn_105_mem);
end

assign tapIn_105 = tapIn_105_mem[d_index];

// Load tapIn_106
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap106.hex",tapIn_106_mem);
end

assign tapIn_106 = tapIn_106_mem[d_index];

// Load tapIn_107
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap107.hex",tapIn_107_mem);
end

assign tapIn_107 = tapIn_107_mem[d_index];

// Load tapIn_108
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap108.hex",tapIn_108_mem);
end

assign tapIn_108 = tapIn_108_mem[d_index];

// Load tapIn_109
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap109.hex",tapIn_109_mem);
end

assign tapIn_109 = tapIn_109_mem[d_index];

// Load tapIn_110
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap110.hex",tapIn_110_mem);
end

assign tapIn_110 = tapIn_110_mem[d_index];

// Load tapIn_111
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap111.hex",tapIn_111_mem);
end

assign tapIn_111 = tapIn_111_mem[d_index];

// Load tapIn_112
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap112.hex",tapIn_112_mem);
end

assign tapIn_112 = tapIn_112_mem[d_index];

// Load tapIn_113
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap113.hex",tapIn_113_mem);
end

assign tapIn_113 = tapIn_113_mem[d_index];

// Load tapIn_114
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap114.hex",tapIn_114_mem);
end

assign tapIn_114 = tapIn_114_mem[d_index];

// Load tapIn_115
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap115.hex",tapIn_115_mem);
end

assign tapIn_115 = tapIn_115_mem[d_index];

// Load tapIn_116
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap116.hex",tapIn_116_mem);
end

assign tapIn_116 = tapIn_116_mem[d_index];

// Load tapIn_117
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap117.hex",tapIn_117_mem);
end

assign tapIn_117 = tapIn_117_mem[d_index];

// Load tapIn_118
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap118.hex",tapIn_118_mem);
end

assign tapIn_118 = tapIn_118_mem[d_index];

// Load tapIn_119
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap119.hex",tapIn_119_mem);
end

assign tapIn_119 = tapIn_119_mem[d_index];

// Load tapIn_120
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap120.hex",tapIn_120_mem);
end

assign tapIn_120 = tapIn_120_mem[d_index];

// Load tapIn_121
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap121.hex",tapIn_121_mem);
end

assign tapIn_121 = tapIn_121_mem[d_index];

// Load tapIn_122
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap122.hex",tapIn_122_mem);
end

assign tapIn_122 = tapIn_122_mem[d_index];

// Load tapIn_123
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap123.hex",tapIn_123_mem);
end

assign tapIn_123 = tapIn_123_mem[d_index];

// Load tapIn_124
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap124.hex",tapIn_124_mem);
end

assign tapIn_124 = tapIn_124_mem[d_index];

// Load tapIn_125
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap125.hex",tapIn_125_mem);
end

assign tapIn_125 = tapIn_125_mem[d_index];

// Load tapIn_126
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap126.hex",tapIn_126_mem);
end

assign tapIn_126 = tapIn_126_mem[d_index];

// Load tapIn_127
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/tap127.hex",tapIn_127_mem);
end

assign tapIn_127 = tapIn_127_mem[d_index];

// Load biasIn_0
initial begin
  $readmemh("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/bias.hex",biasIn_0_mem);
end

assign biasIn_0 = biasIn_0_mem[counter];

// Store Store dataOut_0
initial begin
  rout1_fptr = $fopen("/home/andy/IdeaProjects/NeuralHDL/tests/neuronStage/data/rout1.hex","w");
end

always @(posedge clk) begin
  if (reset) begin
    
  end
  else begin
    $fdisplay(rout1_fptr,"%h ",dataOut_0);
  end
end

// Counter to Index Test
always @(posedge clk) begin
  if (reset) begin
    counter <= 32'd0;
  end
  else begin
    counter <= counter[31:0] + 32'd1;
  end
end

// Initial Statement
initial begin
  
end


// DUT
endmodule

